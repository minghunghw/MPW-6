# Confidential Information of Artisan Components, Inc.
# Use subject to Artisan Components license.
# Copyright (c) 2022 Artisan Components, Inc.

# ACI Version 2008Q3V1

# Reifier 1.1.2

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;

BUSBITCHARS "[]" ;

#name: High Speed/Density Single Port SRAM Generator|IBM CMRF8SF-LPVT Process
#version: 2008Q3V1
#comment: 
#configuration:  -instname RA1SHD -words 4096 -bits 8 -frequency 1 -ring_width 2.0 -mux 16 -write_mask off -wp_size 8 -top_layer met4 -power_type rings -horiz met3 -vert met4 -cust_comment "" -bus_notation on -left_bus_delim "[" -right_bus_delim "]" -pwr_gnd_rename "VDD:VDD,GND:VSS" -prefix "" -pin_space 0.0 -name_case upper -check_instname on -diodes on -inside_ring_type GND -drive 6 -asvm on -corners ff_1p32v_m40c,ff_1p65v_125c,tt_1p2v_25c,ss_1p08v_125c
MACRO RA1SHD
  FOREIGN RA1SHD 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 240.6 BY 517.18 ;
  CLASS RING ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN A[0] ;
    PORT
      LAYER M1 ;
      RECT 137.81 6.24 138.41 6.84 ;
      LAYER M2 ;
      RECT 137.81 6.24 138.41 6.84 ;
      LAYER M3 ;
      RECT 137.81 6.24 138.41 6.84 ;
      LAYER M4 ;
      RECT 137.81 6.24 138.41 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END A[0]
  PIN A[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN A[10] ;
    PORT
      LAYER M4 ;
      RECT 93.61 6.24 94.21 6.84 ;
      LAYER M3 ;
      RECT 93.61 6.24 94.21 6.84 ;
      LAYER M2 ;
      RECT 93.61 6.24 94.21 6.84 ;
      LAYER M1 ;
      RECT 93.61 6.24 94.21 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END A[10]
  PIN A[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN A[11] ;
    PORT
      LAYER M4 ;
      RECT 90.21 6.24 90.81 6.84 ;
      LAYER M3 ;
      RECT 90.21 6.24 90.81 6.84 ;
      LAYER M2 ;
      RECT 90.21 6.24 90.81 6.84 ;
      LAYER M1 ;
      RECT 90.21 6.24 90.81 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END A[11]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN A[1] ;
    PORT
      LAYER M1 ;
      RECT 134.41 6.24 135.01 6.84 ;
      LAYER M2 ;
      RECT 134.41 6.24 135.01 6.84 ;
      LAYER M3 ;
      RECT 134.41 6.24 135.01 6.84 ;
      LAYER M4 ;
      RECT 134.41 6.24 135.01 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN A[2] ;
    PORT
      LAYER M1 ;
      RECT 131.01 6.24 131.61 6.84 ;
      LAYER M2 ;
      RECT 131.01 6.24 131.61 6.84 ;
      LAYER M3 ;
      RECT 131.01 6.24 131.61 6.84 ;
      LAYER M4 ;
      RECT 131.01 6.24 131.61 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN A[3] ;
    PORT
      LAYER M1 ;
      RECT 127.61 6.24 128.21 6.84 ;
      LAYER M2 ;
      RECT 127.61 6.24 128.21 6.84 ;
      LAYER M3 ;
      RECT 127.61 6.24 128.21 6.84 ;
      LAYER M4 ;
      RECT 127.61 6.24 128.21 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN A[4] ;
    PORT
      LAYER M4 ;
      RECT 120.81 6.24 121.41 6.84 ;
      LAYER M3 ;
      RECT 120.81 6.24 121.41 6.84 ;
      LAYER M2 ;
      RECT 120.81 6.24 121.41 6.84 ;
      LAYER M1 ;
      RECT 120.81 6.24 121.41 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN A[5] ;
    PORT
      LAYER M4 ;
      RECT 117.41 6.24 118.01 6.84 ;
      LAYER M3 ;
      RECT 117.41 6.24 118.01 6.84 ;
      LAYER M2 ;
      RECT 117.41 6.24 118.01 6.84 ;
      LAYER M1 ;
      RECT 117.41 6.24 118.01 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN A[6] ;
    PORT
      LAYER M4 ;
      RECT 114.01 6.24 114.61 6.84 ;
      LAYER M3 ;
      RECT 114.01 6.24 114.61 6.84 ;
      LAYER M2 ;
      RECT 114.01 6.24 114.61 6.84 ;
      LAYER M1 ;
      RECT 114.01 6.24 114.61 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN A[7] ;
    PORT
      LAYER M4 ;
      RECT 107.21 6.24 107.81 6.84 ;
      LAYER M3 ;
      RECT 107.21 6.24 107.81 6.84 ;
      LAYER M2 ;
      RECT 107.21 6.24 107.81 6.84 ;
      LAYER M1 ;
      RECT 107.21 6.24 107.81 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN A[8] ;
    PORT
      LAYER M4 ;
      RECT 103.81 6.24 104.41 6.84 ;
      LAYER M3 ;
      RECT 103.81 6.24 104.41 6.84 ;
      LAYER M2 ;
      RECT 103.81 6.24 104.41 6.84 ;
      LAYER M1 ;
      RECT 103.81 6.24 104.41 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN A[9] ;
    PORT
      LAYER M4 ;
      RECT 100.41 6.24 101.01 6.84 ;
      LAYER M3 ;
      RECT 100.41 6.24 101.01 6.84 ;
      LAYER M2 ;
      RECT 100.41 6.24 101.01 6.84 ;
      LAYER M1 ;
      RECT 100.41 6.24 101.01 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END A[9]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN CEN ;
    PORT
      LAYER M1 ;
      RECT 144.01 6.24 144.61 6.84 ;
      LAYER M2 ;
      RECT 144.01 6.24 144.61 6.84 ;
      LAYER M3 ;
      RECT 144.01 6.24 144.61 6.84 ;
      LAYER M4 ;
      RECT 144.01 6.24 144.61 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END CEN
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN CLK ;
    PORT
      LAYER M1 ;
      RECT 152.89 6.24 153.49 6.84 ;
      LAYER M2 ;
      RECT 152.89 6.24 153.49 6.84 ;
      LAYER M3 ;
      RECT 152.89 6.24 153.49 6.84 ;
      LAYER M4 ;
      RECT 152.89 6.24 153.49 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END CLK
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN D[0] ;
    PORT
      LAYER M4 ;
      RECT 23.71 6.24 24.31 6.84 ;
      LAYER M3 ;
      RECT 23.71 6.24 24.31 6.84 ;
      LAYER M2 ;
      RECT 23.71 6.24 24.31 6.84 ;
      LAYER M1 ;
      RECT 23.71 6.24 24.31 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END D[0]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN D[1] ;
    PORT
      LAYER M4 ;
      RECT 30.91 6.24 31.51 6.84 ;
      LAYER M3 ;
      RECT 30.91 6.24 31.51 6.84 ;
      LAYER M2 ;
      RECT 30.91 6.24 31.51 6.84 ;
      LAYER M1 ;
      RECT 30.91 6.24 31.51 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN D[2] ;
    PORT
      LAYER M4 ;
      RECT 63.31 6.24 63.91 6.84 ;
      LAYER M3 ;
      RECT 63.31 6.24 63.91 6.84 ;
      LAYER M2 ;
      RECT 63.31 6.24 63.91 6.84 ;
      LAYER M1 ;
      RECT 63.31 6.24 63.91 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN D[3] ;
    PORT
      LAYER M4 ;
      RECT 70.51 6.24 71.11 6.84 ;
      LAYER M3 ;
      RECT 70.51 6.24 71.11 6.84 ;
      LAYER M2 ;
      RECT 70.51 6.24 71.11 6.84 ;
      LAYER M1 ;
      RECT 70.51 6.24 71.11 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN D[4] ;
    PORT
      LAYER M1 ;
      RECT 169.49 6.24 170.09 6.84 ;
      LAYER M2 ;
      RECT 169.49 6.24 170.09 6.84 ;
      LAYER M3 ;
      RECT 169.49 6.24 170.09 6.84 ;
      LAYER M4 ;
      RECT 169.49 6.24 170.09 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN D[5] ;
    PORT
      LAYER M1 ;
      RECT 176.69 6.24 177.29 6.84 ;
      LAYER M2 ;
      RECT 176.69 6.24 177.29 6.84 ;
      LAYER M3 ;
      RECT 176.69 6.24 177.29 6.84 ;
      LAYER M4 ;
      RECT 176.69 6.24 177.29 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN D[6] ;
    PORT
      LAYER M1 ;
      RECT 209.09 6.24 209.69 6.84 ;
      LAYER M2 ;
      RECT 209.09 6.24 209.69 6.84 ;
      LAYER M3 ;
      RECT 209.09 6.24 209.69 6.84 ;
      LAYER M4 ;
      RECT 209.09 6.24 209.69 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN D[7] ;
    PORT
      LAYER M1 ;
      RECT 216.29 6.24 216.89 6.84 ;
      LAYER M2 ;
      RECT 216.29 6.24 216.89 6.84 ;
      LAYER M3 ;
      RECT 216.29 6.24 216.89 6.84 ;
      LAYER M4 ;
      RECT 216.29 6.24 216.89 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END D[7]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN Q[0] ;
    PORT
      LAYER M4 ;
      RECT 26.11 6.24 26.71 6.84 ;
      LAYER M3 ;
      RECT 26.11 6.24 26.71 6.84 ;
      LAYER M2 ;
      RECT 26.11 6.24 26.71 6.84 ;
      LAYER M1 ;
      RECT 26.11 6.24 26.71 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END Q[0]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN Q[1] ;
    PORT
      LAYER M4 ;
      RECT 28.51 6.24 29.11 6.84 ;
      LAYER M3 ;
      RECT 28.51 6.24 29.11 6.84 ;
      LAYER M2 ;
      RECT 28.51 6.24 29.11 6.84 ;
      LAYER M1 ;
      RECT 28.51 6.24 29.11 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN Q[2] ;
    PORT
      LAYER M4 ;
      RECT 65.71 6.24 66.31 6.84 ;
      LAYER M3 ;
      RECT 65.71 6.24 66.31 6.84 ;
      LAYER M2 ;
      RECT 65.71 6.24 66.31 6.84 ;
      LAYER M1 ;
      RECT 65.71 6.24 66.31 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN Q[3] ;
    PORT
      LAYER M4 ;
      RECT 68.11 6.24 68.71 6.84 ;
      LAYER M3 ;
      RECT 68.11 6.24 68.71 6.84 ;
      LAYER M2 ;
      RECT 68.11 6.24 68.71 6.84 ;
      LAYER M1 ;
      RECT 68.11 6.24 68.71 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN Q[4] ;
    PORT
      LAYER M1 ;
      RECT 171.89 6.24 172.49 6.84 ;
      LAYER M2 ;
      RECT 171.89 6.24 172.49 6.84 ;
      LAYER M3 ;
      RECT 171.89 6.24 172.49 6.84 ;
      LAYER M4 ;
      RECT 171.89 6.24 172.49 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN Q[5] ;
    PORT
      LAYER M1 ;
      RECT 174.29 6.24 174.89 6.84 ;
      LAYER M2 ;
      RECT 174.29 6.24 174.89 6.84 ;
      LAYER M3 ;
      RECT 174.29 6.24 174.89 6.84 ;
      LAYER M4 ;
      RECT 174.29 6.24 174.89 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN Q[6] ;
    PORT
      LAYER M1 ;
      RECT 211.49 6.24 212.09 6.84 ;
      LAYER M2 ;
      RECT 211.49 6.24 212.09 6.84 ;
      LAYER M3 ;
      RECT 211.49 6.24 212.09 6.84 ;
      LAYER M4 ;
      RECT 211.49 6.24 212.09 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN Q[7] ;
    PORT
      LAYER M1 ;
      RECT 213.89 6.24 214.49 6.84 ;
      LAYER M2 ;
      RECT 213.89 6.24 214.49 6.84 ;
      LAYER M3 ;
      RECT 213.89 6.24 214.49 6.84 ;
      LAYER M4 ;
      RECT 213.89 6.24 214.49 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END Q[7]
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    FOREIGN WEN ;
    PORT
      LAYER M1 ;
      RECT 149.27 6.24 149.87 6.84 ;
      LAYER M2 ;
      RECT 149.27 6.24 149.87 6.84 ;
      LAYER M3 ;
      RECT 149.27 6.24 149.87 6.84 ;
      LAYER M4 ;
      RECT 149.27 6.24 149.87 6.84 ;
      END
    ANTENNAGATEAREA 0.0384 ;
    ANTENNADIFFAREA 0.0784 ;
    END WEN
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER M3 ;
      RECT 3.12 512.06 237.48 514.06 ;
      END
    PORT
      LAYER M3 ;
      RECT 3.12 3.12 237.48 5.12 ;
      END
    PORT
      LAYER M4 ;
      RECT 235.48 3.12 237.48 514.06 ;
      END
    PORT
      LAYER M4 ;
      RECT 3.12 3.12 5.12 514.06 ;
      END
    END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER M3 ;
      RECT 0.0 515.18 240.6 517.18 ;
      END
    PORT
      LAYER M3 ;
      RECT 0.0 0.0 240.6 2.0 ;
      END
    PORT
      LAYER M4 ;
      RECT 238.6 0.0 240.6 517.18 ;
      END
    PORT
      LAYER M4 ;
      RECT 0.0 0.0 2.0 517.18 ;
      END
    END VDD
  OBS
    #core
    LAYER V1 ;
    RECT 6.24 6.24 234.36 510.94 ;
    LAYER V2 ;
    RECT 6.24 6.24 234.36 510.94 ;
    LAYER V3 ;
    RECT 6.24 6.24 234.36 510.94 ;
    LAYER OVERLAP ;
    RECT 6.24 6.24 234.36 510.94 ;
    #notched core
    LAYER M1 SPACING 0.16 ;
    POLYGON 6.24 510.94 6.24 6.24 23.55 6.24 23.55 7.0 24.47 7.0 24.47 6.24
      25.95 6.24 25.95 7.0 26.87 7.0 26.87 6.24 28.35 6.24 28.35 7.0
      29.27 7.0 29.27 6.24 30.75 6.24 30.75 7.0 31.67 7.0 31.67 6.24
      63.15 6.24 63.15 7.0 64.07 7.0 64.07 6.24 65.55 6.24 65.55 7.0
      66.47 7.0 66.47 6.24 67.95 6.24 67.95 7.0 68.87 7.0 68.87 6.24
      70.35 6.24 70.35 7.0 71.27 7.0 71.27 6.24 90.05 6.24 90.05 7.0
      90.97 7.0 90.97 6.24 93.45 6.24 93.45 7.0 94.37 7.0 94.37 6.24
      100.25 6.24 100.25 7.0 101.17 7.0 101.17 6.24 103.65 6.24 103.65 7.0
      104.57 7.0 104.57 6.24 107.05 6.24 107.05 7.0 107.97 7.0 107.97 6.24
      113.85 6.24 113.85 7.0 114.77 7.0 114.77 6.24 117.25 6.24 117.25 7.0
      118.17 7.0 118.17 6.24 120.65 6.24 120.65 7.0 121.57 7.0 121.57 6.24
      127.45 6.24 127.45 7.0 128.37 7.0 128.37 6.24 130.85 6.24 130.85 7.0
      131.77 7.0 131.77 6.24 134.25 6.24 134.25 7.0 135.17 7.0 135.17 6.24
      137.65 6.24 137.65 7.0 138.57 7.0 138.57 6.24 143.85 6.24 143.85 7.0
      144.77 7.0 144.77 6.24 149.11 6.24 149.11 7.0 150.03 7.0 150.03 6.24
      152.73 6.24 152.73 7.0 153.65 7.0 153.65 6.24 169.33 6.24 169.33 7.0
      170.25 7.0 170.25 6.24 171.73 6.24 171.73 7.0 172.65 7.0 172.65 6.24
      174.13 6.24 174.13 7.0 175.05 7.0 175.05 6.24 176.53 6.24 176.53 7.0
      177.45 7.0 177.45 6.24 208.93 6.24 208.93 7.0 209.85 7.0 209.85 6.24
      211.33 6.24 211.33 7.0 212.25 7.0 212.25 6.24 213.73 6.24 213.73 7.0
      214.65 7.0 214.65 6.24 216.13 6.24 216.13 7.0 217.05 7.0 217.05 6.24
      234.36 6.24 234.36 510.94 ;
    #notched core
    LAYER M2 SPACING 0.2 ;
    POLYGON 6.24 510.94 6.24 6.24 23.51 6.24 23.51 7.04 24.51 7.04 24.51 6.24
      25.91 6.24 25.91 7.04 26.91 7.04 26.91 6.24 28.31 6.24 28.31 7.04
      29.31 7.04 29.31 6.24 30.71 6.24 30.71 7.04 31.71 7.04 31.71 6.24
      63.11 6.24 63.11 7.04 64.11 7.04 64.11 6.24 65.51 6.24 65.51 7.04
      66.51 7.04 66.51 6.24 67.91 6.24 67.91 7.04 68.91 7.04 68.91 6.24
      70.31 6.24 70.31 7.04 71.31 7.04 71.31 6.24 90.01 6.24 90.01 7.04
      91.01 7.04 91.01 6.24 93.41 6.24 93.41 7.04 94.41 7.04 94.41 6.24
      100.21 6.24 100.21 7.04 101.21 7.04 101.21 6.24 103.61 6.24 103.61 7.04
      104.61 7.04 104.61 6.24 107.01 6.24 107.01 7.04 108.01 7.04 108.01 6.24
      113.81 6.24 113.81 7.04 114.81 7.04 114.81 6.24 117.21 6.24 117.21 7.04
      118.21 7.04 118.21 6.24 120.61 6.24 120.61 7.04 121.61 7.04 121.61 6.24
      127.41 6.24 127.41 7.04 128.41 7.04 128.41 6.24 130.81 6.24 130.81 7.04
      131.81 7.04 131.81 6.24 134.21 6.24 134.21 7.04 135.21 7.04 135.21 6.24
      137.61 6.24 137.61 7.04 138.61 7.04 138.61 6.24 143.81 6.24 143.81 7.04
      144.81 7.04 144.81 6.24 149.07 6.24 149.07 7.04 150.07 7.04 150.07 6.24
      152.69 6.24 152.69 7.04 153.69 7.04 153.69 6.24 169.29 6.24 169.29 7.04
      170.29 7.04 170.29 6.24 171.69 6.24 171.69 7.04 172.69 7.04 172.69 6.24
      174.09 6.24 174.09 7.04 175.09 7.04 175.09 6.24 176.49 6.24 176.49 7.04
      177.49 7.04 177.49 6.24 208.89 6.24 208.89 7.04 209.89 7.04 209.89 6.24
      211.29 6.24 211.29 7.04 212.29 7.04 212.29 6.24 213.69 6.24 213.69 7.04
      214.69 7.04 214.69 6.24 216.09 6.24 216.09 7.04 217.09 7.04 217.09 6.24
      234.36 6.24 234.36 510.94 ;
    #notched core
    LAYER M3 SPACING 0.2 ;
    POLYGON 6.24 510.94 6.24 6.24 23.51 6.24 23.51 7.04 24.51 7.04 24.51 6.24
      25.91 6.24 25.91 7.04 26.91 7.04 26.91 6.24 28.31 6.24 28.31 7.04
      29.31 7.04 29.31 6.24 30.71 6.24 30.71 7.04 31.71 7.04 31.71 6.24
      63.11 6.24 63.11 7.04 64.11 7.04 64.11 6.24 65.51 6.24 65.51 7.04
      66.51 7.04 66.51 6.24 67.91 6.24 67.91 7.04 68.91 7.04 68.91 6.24
      70.31 6.24 70.31 7.04 71.31 7.04 71.31 6.24 90.01 6.24 90.01 7.04
      91.01 7.04 91.01 6.24 93.41 6.24 93.41 7.04 94.41 7.04 94.41 6.24
      100.21 6.24 100.21 7.04 101.21 7.04 101.21 6.24 103.61 6.24 103.61 7.04
      104.61 7.04 104.61 6.24 107.01 6.24 107.01 7.04 108.01 7.04 108.01 6.24
      113.81 6.24 113.81 7.04 114.81 7.04 114.81 6.24 117.21 6.24 117.21 7.04
      118.21 7.04 118.21 6.24 120.61 6.24 120.61 7.04 121.61 7.04 121.61 6.24
      127.41 6.24 127.41 7.04 128.41 7.04 128.41 6.24 130.81 6.24 130.81 7.04
      131.81 7.04 131.81 6.24 134.21 6.24 134.21 7.04 135.21 7.04 135.21 6.24
      137.61 6.24 137.61 7.04 138.61 7.04 138.61 6.24 143.81 6.24 143.81 7.04
      144.81 7.04 144.81 6.24 149.07 6.24 149.07 7.04 150.07 7.04 150.07 6.24
      152.69 6.24 152.69 7.04 153.69 7.04 153.69 6.24 169.29 6.24 169.29 7.04
      170.29 7.04 170.29 6.24 171.69 6.24 171.69 7.04 172.69 7.04 172.69 6.24
      174.09 6.24 174.09 7.04 175.09 7.04 175.09 6.24 176.49 6.24 176.49 7.04
      177.49 7.04 177.49 6.24 208.89 6.24 208.89 7.04 209.89 7.04 209.89 6.24
      211.29 6.24 211.29 7.04 212.29 7.04 212.29 6.24 213.69 6.24 213.69 7.04
      214.69 7.04 214.69 6.24 216.09 6.24 216.09 7.04 217.09 7.04 217.09 6.24
      234.36 6.24 234.36 510.94 ;
    #notched core
    LAYER M4 SPACING 0.2 ;
    POLYGON 6.24 510.94 6.24 6.24 23.51 6.24 23.51 7.04 24.51 7.04 24.51 6.24
      25.91 6.24 25.91 7.04 26.91 7.04 26.91 6.24 28.31 6.24 28.31 7.04
      29.31 7.04 29.31 6.24 30.71 6.24 30.71 7.04 31.71 7.04 31.71 6.24
      63.11 6.24 63.11 7.04 64.11 7.04 64.11 6.24 65.51 6.24 65.51 7.04
      66.51 7.04 66.51 6.24 67.91 6.24 67.91 7.04 68.91 7.04 68.91 6.24
      70.31 6.24 70.31 7.04 71.31 7.04 71.31 6.24 90.01 6.24 90.01 7.04
      91.01 7.04 91.01 6.24 93.41 6.24 93.41 7.04 94.41 7.04 94.41 6.24
      100.21 6.24 100.21 7.04 101.21 7.04 101.21 6.24 103.61 6.24 103.61 7.04
      104.61 7.04 104.61 6.24 107.01 6.24 107.01 7.04 108.01 7.04 108.01 6.24
      113.81 6.24 113.81 7.04 114.81 7.04 114.81 6.24 117.21 6.24 117.21 7.04
      118.21 7.04 118.21 6.24 120.61 6.24 120.61 7.04 121.61 7.04 121.61 6.24
      127.41 6.24 127.41 7.04 128.41 7.04 128.41 6.24 130.81 6.24 130.81 7.04
      131.81 7.04 131.81 6.24 134.21 6.24 134.21 7.04 135.21 7.04 135.21 6.24
      137.61 6.24 137.61 7.04 138.61 7.04 138.61 6.24 143.81 6.24 143.81 7.04
      144.81 7.04 144.81 6.24 149.07 6.24 149.07 7.04 150.07 7.04 150.07 6.24
      152.69 6.24 152.69 7.04 153.69 7.04 153.69 6.24 169.29 6.24 169.29 7.04
      170.29 7.04 170.29 6.24 171.69 6.24 171.69 7.04 172.69 7.04 172.69 6.24
      174.09 6.24 174.09 7.04 175.09 7.04 175.09 6.24 176.49 6.24 176.49 7.04
      177.49 7.04 177.49 6.24 208.89 6.24 208.89 7.04 209.89 7.04 209.89 6.24
      211.29 6.24 211.29 7.04 212.29 7.04 212.29 6.24 213.69 6.24 213.69 7.04
      214.69 7.04 214.69 6.24 216.09 6.24 216.09 7.04 217.09 7.04 217.09 6.24
      234.36 6.24 234.36 510.94 ;
    #power fingers
    LAYER M4 ;
    RECT 9.81 510.94 11.81 517.18 ;
    LAYER M4 ;
    RECT 14.61 510.94 16.61 517.18 ;
    LAYER M4 ;
    RECT 19.41 510.94 21.41 517.18 ;
    LAYER M4 ;
    RECT 24.21 510.94 26.21 517.18 ;
    LAYER M4 ;
    RECT 29.01 510.94 31.01 517.18 ;
    LAYER M4 ;
    RECT 33.81 510.94 35.81 517.18 ;
    LAYER M4 ;
    RECT 38.61 510.94 40.61 517.18 ;
    LAYER M4 ;
    RECT 43.41 510.94 45.41 517.18 ;
    LAYER M4 ;
    RECT 49.41 510.94 51.41 517.18 ;
    LAYER M4 ;
    RECT 54.21 510.94 56.21 517.18 ;
    LAYER M4 ;
    RECT 59.01 510.94 61.01 517.18 ;
    LAYER M4 ;
    RECT 63.81 510.94 65.81 517.18 ;
    LAYER M4 ;
    RECT 68.61 510.94 70.61 517.18 ;
    LAYER M4 ;
    RECT 73.41 510.94 75.41 517.18 ;
    LAYER M4 ;
    RECT 78.21 510.94 80.21 517.18 ;
    LAYER M4 ;
    RECT 83.01 510.94 85.01 517.18 ;
    LAYER M4 ;
    RECT 87.81 510.94 88.61 517.18 ;
    LAYER M4 ;
    RECT 90.81 510.94 91.91 517.18 ;
    LAYER M4 ;
    RECT 94.21 510.94 95.31 517.18 ;
    LAYER M4 ;
    RECT 97.61 510.94 98.71 517.18 ;
    LAYER M4 ;
    RECT 101.01 510.94 102.11 517.18 ;
    LAYER M4 ;
    RECT 104.41 510.94 105.51 517.18 ;
    LAYER M4 ;
    RECT 107.81 510.94 108.91 517.18 ;
    LAYER M4 ;
    RECT 111.21 510.94 114.01 517.18 ;
    LAYER M4 ;
    RECT 118.01 510.94 120.81 517.18 ;
    LAYER M4 ;
    RECT 124.81 510.94 127.61 517.18 ;
    LAYER M4 ;
    RECT 131.61 510.94 134.41 517.18 ;
    LAYER M4 ;
    RECT 138.41 510.94 141.65 517.18 ;
    LAYER M4 ;
    RECT 144.17 510.94 145.49 517.18 ;
    LAYER M4 ;
    RECT 148.01 510.94 149.33 517.18 ;
    LAYER M4 ;
    RECT 151.99 510.94 152.79 517.18 ;
    LAYER M4 ;
    RECT 155.59 510.94 157.59 517.18 ;
    LAYER M4 ;
    RECT 160.39 510.94 162.39 517.18 ;
    LAYER M4 ;
    RECT 165.19 510.94 167.19 517.18 ;
    LAYER M4 ;
    RECT 169.99 510.94 171.99 517.18 ;
    LAYER M4 ;
    RECT 174.79 510.94 176.79 517.18 ;
    LAYER M4 ;
    RECT 179.59 510.94 181.59 517.18 ;
    LAYER M4 ;
    RECT 184.39 510.94 186.39 517.18 ;
    LAYER M4 ;
    RECT 189.19 510.94 191.19 517.18 ;
    LAYER M4 ;
    RECT 195.19 510.94 197.19 517.18 ;
    LAYER M4 ;
    RECT 199.99 510.94 201.99 517.18 ;
    LAYER M4 ;
    RECT 204.79 510.94 206.79 517.18 ;
    LAYER M4 ;
    RECT 209.59 510.94 211.59 517.18 ;
    LAYER M4 ;
    RECT 214.39 510.94 216.39 517.18 ;
    LAYER M4 ;
    RECT 219.19 510.94 221.19 517.18 ;
    LAYER M4 ;
    RECT 223.99 510.94 225.99 517.18 ;
    LAYER M4 ;
    RECT 228.79 510.94 230.79 517.18 ;
    LAYER M4 ;
    RECT 9.81 0.0 11.79 6.24 ;
    LAYER M4 ;
    RECT 14.61 0.0 16.59 6.24 ;
    LAYER M4 ;
    RECT 19.81 0.0 21.41 6.24 ;
    LAYER M4 ;
    RECT 24.71 0.0 25.71 6.24 ;
    LAYER M4 ;
    RECT 29.51 0.0 30.51 6.24 ;
    LAYER M4 ;
    RECT 33.84 0.0 35.81 6.24 ;
    LAYER M4 ;
    RECT 38.63 0.0 40.61 6.24 ;
    LAYER M4 ;
    RECT 43.43 0.0 45.41 6.24 ;
    LAYER M4 ;
    RECT 49.41 0.0 51.39 6.24 ;
    LAYER M4 ;
    RECT 54.21 0.0 56.19 6.24 ;
    LAYER M4 ;
    RECT 59.01 0.0 60.98 6.24 ;
    LAYER M4 ;
    RECT 64.31 0.0 65.31 6.24 ;
    LAYER M4 ;
    RECT 69.11 0.0 70.11 6.24 ;
    LAYER M4 ;
    RECT 73.44 0.0 75.41 6.24 ;
    LAYER M4 ;
    RECT 78.23 0.0 80.21 6.24 ;
    LAYER M4 ;
    RECT 83.03 0.0 85.01 6.24 ;
    LAYER M4 ;
    RECT 87.21 0.0 88.01 6.24 ;
    LAYER M4 ;
    RECT 91.23 0.0 93.19 6.24 ;
    LAYER M4 ;
    RECT 98.01 0.0 99.99 6.24 ;
    LAYER M4 ;
    RECT 104.83 0.0 106.79 6.24 ;
    LAYER M4 ;
    RECT 111.61 0.0 113.59 6.24 ;
    LAYER M4 ;
    RECT 118.43 0.0 120.39 6.24 ;
    LAYER M4 ;
    RECT 125.21 0.0 127.19 6.24 ;
    LAYER M4 ;
    RECT 132.03 0.0 133.99 6.24 ;
    LAYER M4 ;
    RECT 138.83 0.0 140.83 6.24 ;
    LAYER M4 ;
    RECT 145.01 0.0 145.61 6.24 ;
    LAYER M4 ;
    RECT 148.01 0.0 148.87 6.24 ;
    LAYER M4 ;
    RECT 155.59 0.0 157.57 6.24 ;
    LAYER M4 ;
    RECT 160.39 0.0 162.37 6.24 ;
    LAYER M4 ;
    RECT 165.19 0.0 167.16 6.24 ;
    LAYER M4 ;
    RECT 170.49 0.0 171.49 6.24 ;
    LAYER M4 ;
    RECT 175.29 0.0 176.29 6.24 ;
    LAYER M4 ;
    RECT 179.62 0.0 181.59 6.24 ;
    LAYER M4 ;
    RECT 184.41 0.0 186.39 6.24 ;
    LAYER M4 ;
    RECT 189.21 0.0 191.19 6.24 ;
    LAYER M4 ;
    RECT 195.19 0.0 197.17 6.24 ;
    LAYER M4 ;
    RECT 199.99 0.0 201.97 6.24 ;
    LAYER M4 ;
    RECT 204.79 0.0 206.76 6.24 ;
    LAYER M4 ;
    RECT 210.09 0.0 211.09 6.24 ;
    LAYER M4 ;
    RECT 214.89 0.0 215.89 6.24 ;
    LAYER M4 ;
    RECT 219.21 0.0 221.19 6.24 ;
    LAYER M4 ;
    RECT 224.01 0.0 225.99 6.24 ;
    LAYER M4 ;
    RECT 228.81 0.0 230.79 6.24 ;
    LAYER M3 ;
    RECT 234.36 7.94 240.6 9.14 ;
    LAYER M3 ;
    RECT 234.36 17.26 240.6 18.46 ;
    LAYER M3 ;
    RECT 234.36 25.81 240.6 27.81 ;
    LAYER M3 ;
    RECT 234.36 35.91 240.6 36.91 ;
    LAYER M3 ;
    RECT 234.36 50.24 240.6 51.24 ;
    LAYER M3 ;
    RECT 234.36 57.02 240.6 58.02 ;
    LAYER M3 ;
    RECT 234.36 60.6 240.6 61.6 ;
    LAYER M3 ;
    RECT 234.36 62.45 240.6 63.45 ;
    LAYER M3 ;
    RECT 234.36 69.16 240.6 69.96 ;
    LAYER M3 ;
    RECT 234.36 72.56 240.6 73.36 ;
    LAYER M3 ;
    RECT 234.36 75.96 240.6 76.76 ;
    LAYER M3 ;
    RECT 234.36 79.36 240.6 80.16 ;
    LAYER M3 ;
    RECT 234.36 82.76 240.6 83.56 ;
    LAYER M3 ;
    RECT 234.36 86.16 240.6 86.96 ;
    LAYER M3 ;
    RECT 234.36 89.56 240.6 90.36 ;
    LAYER M3 ;
    RECT 234.36 92.96 240.6 93.76 ;
    LAYER M3 ;
    RECT 234.36 96.36 240.6 97.16 ;
    LAYER M3 ;
    RECT 234.36 99.76 240.6 100.56 ;
    LAYER M3 ;
    RECT 234.36 103.16 240.6 103.96 ;
    LAYER M3 ;
    RECT 234.36 106.56 240.6 107.36 ;
    LAYER M3 ;
    RECT 234.36 109.96 240.6 110.76 ;
    LAYER M3 ;
    RECT 234.36 113.36 240.6 114.16 ;
    LAYER M3 ;
    RECT 234.36 116.76 240.6 117.56 ;
    LAYER M3 ;
    RECT 234.36 120.16 240.6 120.96 ;
    LAYER M3 ;
    RECT 234.36 123.56 240.6 124.36 ;
    LAYER M3 ;
    RECT 234.36 126.96 240.6 127.76 ;
    LAYER M3 ;
    RECT 234.36 130.36 240.6 131.16 ;
    LAYER M3 ;
    RECT 234.36 133.76 240.6 134.56 ;
    LAYER M3 ;
    RECT 234.36 137.16 240.6 137.96 ;
    LAYER M3 ;
    RECT 234.36 140.56 240.6 141.36 ;
    LAYER M3 ;
    RECT 234.36 143.96 240.6 144.76 ;
    LAYER M3 ;
    RECT 234.36 147.36 240.6 148.16 ;
    LAYER M3 ;
    RECT 234.36 150.76 240.6 151.56 ;
    LAYER M3 ;
    RECT 234.36 154.16 240.6 154.96 ;
    LAYER M3 ;
    RECT 234.36 157.56 240.6 158.36 ;
    LAYER M3 ;
    RECT 234.36 160.96 240.6 161.76 ;
    LAYER M3 ;
    RECT 234.36 164.36 240.6 165.16 ;
    LAYER M3 ;
    RECT 234.36 167.76 240.6 168.56 ;
    LAYER M3 ;
    RECT 234.36 171.16 240.6 171.96 ;
    LAYER M3 ;
    RECT 234.36 174.56 240.6 175.36 ;
    LAYER M3 ;
    RECT 234.36 177.96 240.6 178.76 ;
    LAYER M3 ;
    RECT 234.36 181.36 240.6 182.16 ;
    LAYER M3 ;
    RECT 234.36 184.76 240.6 185.56 ;
    LAYER M3 ;
    RECT 234.36 188.16 240.6 188.96 ;
    LAYER M3 ;
    RECT 234.36 191.56 240.6 192.36 ;
    LAYER M3 ;
    RECT 234.36 194.96 240.6 195.76 ;
    LAYER M3 ;
    RECT 234.36 198.36 240.6 199.16 ;
    LAYER M3 ;
    RECT 234.36 201.76 240.6 202.56 ;
    LAYER M3 ;
    RECT 234.36 205.16 240.6 205.96 ;
    LAYER M3 ;
    RECT 234.36 208.56 240.6 209.36 ;
    LAYER M3 ;
    RECT 234.36 211.96 240.6 212.76 ;
    LAYER M3 ;
    RECT 234.36 215.36 240.6 216.16 ;
    LAYER M3 ;
    RECT 234.36 218.76 240.6 219.56 ;
    LAYER M3 ;
    RECT 234.36 222.16 240.6 222.96 ;
    LAYER M3 ;
    RECT 234.36 225.56 240.6 226.36 ;
    LAYER M3 ;
    RECT 234.36 228.96 240.6 229.76 ;
    LAYER M3 ;
    RECT 234.36 232.36 240.6 233.16 ;
    LAYER M3 ;
    RECT 234.36 235.76 240.6 236.56 ;
    LAYER M3 ;
    RECT 234.36 239.16 240.6 239.96 ;
    LAYER M3 ;
    RECT 234.36 242.56 240.6 243.36 ;
    LAYER M3 ;
    RECT 234.36 245.96 240.6 246.76 ;
    LAYER M3 ;
    RECT 234.36 249.36 240.6 250.16 ;
    LAYER M3 ;
    RECT 234.36 252.76 240.6 253.56 ;
    LAYER M3 ;
    RECT 234.36 256.16 240.6 256.96 ;
    LAYER M3 ;
    RECT 234.36 259.56 240.6 260.36 ;
    LAYER M3 ;
    RECT 234.36 262.96 240.6 263.76 ;
    LAYER M3 ;
    RECT 234.36 266.36 240.6 267.16 ;
    LAYER M3 ;
    RECT 234.36 269.76 240.6 270.56 ;
    LAYER M3 ;
    RECT 234.36 273.16 240.6 273.96 ;
    LAYER M3 ;
    RECT 234.36 276.56 240.6 277.36 ;
    LAYER M3 ;
    RECT 234.36 279.96 240.6 280.76 ;
    LAYER M3 ;
    RECT 234.36 283.36 240.6 284.16 ;
    LAYER M3 ;
    RECT 234.36 286.76 240.6 287.56 ;
    LAYER M3 ;
    RECT 234.36 290.16 240.6 290.96 ;
    LAYER M3 ;
    RECT 234.36 293.56 240.6 294.36 ;
    LAYER M3 ;
    RECT 234.36 296.96 240.6 297.76 ;
    LAYER M3 ;
    RECT 234.36 300.36 240.6 301.16 ;
    LAYER M3 ;
    RECT 234.36 303.76 240.6 304.56 ;
    LAYER M3 ;
    RECT 234.36 307.16 240.6 307.96 ;
    LAYER M3 ;
    RECT 234.36 310.56 240.6 311.36 ;
    LAYER M3 ;
    RECT 234.36 313.96 240.6 314.76 ;
    LAYER M3 ;
    RECT 234.36 317.36 240.6 318.16 ;
    LAYER M3 ;
    RECT 234.36 320.76 240.6 321.56 ;
    LAYER M3 ;
    RECT 234.36 324.16 240.6 324.96 ;
    LAYER M3 ;
    RECT 234.36 327.56 240.6 328.36 ;
    LAYER M3 ;
    RECT 234.36 330.96 240.6 331.76 ;
    LAYER M3 ;
    RECT 234.36 334.36 240.6 335.16 ;
    LAYER M3 ;
    RECT 234.36 337.76 240.6 338.56 ;
    LAYER M3 ;
    RECT 234.36 341.16 240.6 341.96 ;
    LAYER M3 ;
    RECT 234.36 344.56 240.6 345.36 ;
    LAYER M3 ;
    RECT 234.36 347.96 240.6 348.76 ;
    LAYER M3 ;
    RECT 234.36 351.36 240.6 352.16 ;
    LAYER M3 ;
    RECT 234.36 354.76 240.6 355.56 ;
    LAYER M3 ;
    RECT 234.36 358.16 240.6 358.96 ;
    LAYER M3 ;
    RECT 234.36 361.56 240.6 362.36 ;
    LAYER M3 ;
    RECT 234.36 364.96 240.6 365.76 ;
    LAYER M3 ;
    RECT 234.36 368.36 240.6 369.16 ;
    LAYER M3 ;
    RECT 234.36 371.76 240.6 372.56 ;
    LAYER M3 ;
    RECT 234.36 375.16 240.6 375.96 ;
    LAYER M3 ;
    RECT 234.36 378.56 240.6 379.36 ;
    LAYER M3 ;
    RECT 234.36 381.96 240.6 382.76 ;
    LAYER M3 ;
    RECT 234.36 385.36 240.6 386.16 ;
    LAYER M3 ;
    RECT 234.36 388.76 240.6 389.56 ;
    LAYER M3 ;
    RECT 234.36 392.16 240.6 392.96 ;
    LAYER M3 ;
    RECT 234.36 395.56 240.6 396.36 ;
    LAYER M3 ;
    RECT 234.36 398.96 240.6 399.76 ;
    LAYER M3 ;
    RECT 234.36 402.36 240.6 403.16 ;
    LAYER M3 ;
    RECT 234.36 405.76 240.6 406.56 ;
    LAYER M3 ;
    RECT 234.36 409.16 240.6 409.96 ;
    LAYER M3 ;
    RECT 234.36 412.56 240.6 413.36 ;
    LAYER M3 ;
    RECT 234.36 415.96 240.6 416.76 ;
    LAYER M3 ;
    RECT 234.36 419.36 240.6 420.16 ;
    LAYER M3 ;
    RECT 234.36 422.76 240.6 423.56 ;
    LAYER M3 ;
    RECT 234.36 426.16 240.6 426.96 ;
    LAYER M3 ;
    RECT 234.36 429.56 240.6 430.36 ;
    LAYER M3 ;
    RECT 234.36 432.96 240.6 433.76 ;
    LAYER M3 ;
    RECT 234.36 436.36 240.6 437.16 ;
    LAYER M3 ;
    RECT 234.36 439.76 240.6 440.56 ;
    LAYER M3 ;
    RECT 234.36 443.16 240.6 443.96 ;
    LAYER M3 ;
    RECT 234.36 446.56 240.6 447.36 ;
    LAYER M3 ;
    RECT 234.36 449.96 240.6 450.76 ;
    LAYER M3 ;
    RECT 234.36 453.36 240.6 454.16 ;
    LAYER M3 ;
    RECT 234.36 456.76 240.6 457.56 ;
    LAYER M3 ;
    RECT 234.36 460.16 240.6 460.96 ;
    LAYER M3 ;
    RECT 234.36 463.56 240.6 464.36 ;
    LAYER M3 ;
    RECT 234.36 466.96 240.6 467.76 ;
    LAYER M3 ;
    RECT 234.36 470.36 240.6 471.16 ;
    LAYER M3 ;
    RECT 234.36 473.76 240.6 474.56 ;
    LAYER M3 ;
    RECT 234.36 477.16 240.6 477.96 ;
    LAYER M3 ;
    RECT 234.36 480.56 240.6 481.36 ;
    LAYER M3 ;
    RECT 234.36 483.96 240.6 484.76 ;
    LAYER M3 ;
    RECT 234.36 487.36 240.6 488.16 ;
    LAYER M3 ;
    RECT 234.36 490.76 240.6 491.56 ;
    LAYER M3 ;
    RECT 234.36 494.16 240.6 494.96 ;
    LAYER M3 ;
    RECT 234.36 497.56 240.6 498.36 ;
    LAYER M3 ;
    RECT 234.36 500.96 240.6 501.76 ;
    LAYER M3 ;
    RECT 234.36 504.36 240.6 505.16 ;
    LAYER M3 ;
    RECT 234.36 505.6 240.6 506.0 ;
    LAYER M3 ;
    RECT 234.36 509.0 240.6 509.8 ;
    LAYER M3 ;
    RECT 0.0 7.94 6.24 9.14 ;
    LAYER M3 ;
    RECT 0.0 17.26 6.24 18.46 ;
    LAYER M3 ;
    RECT 0.0 25.81 6.24 27.81 ;
    LAYER M3 ;
    RECT 0.0 35.91 6.24 36.91 ;
    LAYER M3 ;
    RECT 0.0 50.24 6.24 51.24 ;
    LAYER M3 ;
    RECT 0.0 57.02 6.24 58.02 ;
    LAYER M3 ;
    RECT 0.0 60.6 6.24 61.6 ;
    LAYER M3 ;
    RECT 0.0 62.45 6.24 63.45 ;
    LAYER M3 ;
    RECT 0.0 69.16 6.24 69.96 ;
    LAYER M3 ;
    RECT 0.0 72.56 6.24 73.36 ;
    LAYER M3 ;
    RECT 0.0 75.96 6.24 76.76 ;
    LAYER M3 ;
    RECT 0.0 79.36 6.24 80.16 ;
    LAYER M3 ;
    RECT 0.0 82.76 6.24 83.56 ;
    LAYER M3 ;
    RECT 0.0 86.16 6.24 86.96 ;
    LAYER M3 ;
    RECT 0.0 89.56 6.24 90.36 ;
    LAYER M3 ;
    RECT 0.0 92.96 6.24 93.76 ;
    LAYER M3 ;
    RECT 0.0 96.36 6.24 97.16 ;
    LAYER M3 ;
    RECT 0.0 99.76 6.24 100.56 ;
    LAYER M3 ;
    RECT 0.0 103.16 6.24 103.96 ;
    LAYER M3 ;
    RECT 0.0 106.56 6.24 107.36 ;
    LAYER M3 ;
    RECT 0.0 109.96 6.24 110.76 ;
    LAYER M3 ;
    RECT 0.0 113.36 6.24 114.16 ;
    LAYER M3 ;
    RECT 0.0 116.76 6.24 117.56 ;
    LAYER M3 ;
    RECT 0.0 120.16 6.24 120.96 ;
    LAYER M3 ;
    RECT 0.0 123.56 6.24 124.36 ;
    LAYER M3 ;
    RECT 0.0 126.96 6.24 127.76 ;
    LAYER M3 ;
    RECT 0.0 130.36 6.24 131.16 ;
    LAYER M3 ;
    RECT 0.0 133.76 6.24 134.56 ;
    LAYER M3 ;
    RECT 0.0 137.16 6.24 137.96 ;
    LAYER M3 ;
    RECT 0.0 140.56 6.24 141.36 ;
    LAYER M3 ;
    RECT 0.0 143.96 6.24 144.76 ;
    LAYER M3 ;
    RECT 0.0 147.36 6.24 148.16 ;
    LAYER M3 ;
    RECT 0.0 150.76 6.24 151.56 ;
    LAYER M3 ;
    RECT 0.0 154.16 6.24 154.96 ;
    LAYER M3 ;
    RECT 0.0 157.56 6.24 158.36 ;
    LAYER M3 ;
    RECT 0.0 160.96 6.24 161.76 ;
    LAYER M3 ;
    RECT 0.0 164.36 6.24 165.16 ;
    LAYER M3 ;
    RECT 0.0 167.76 6.24 168.56 ;
    LAYER M3 ;
    RECT 0.0 171.16 6.24 171.96 ;
    LAYER M3 ;
    RECT 0.0 174.56 6.24 175.36 ;
    LAYER M3 ;
    RECT 0.0 177.96 6.24 178.76 ;
    LAYER M3 ;
    RECT 0.0 181.36 6.24 182.16 ;
    LAYER M3 ;
    RECT 0.0 184.76 6.24 185.56 ;
    LAYER M3 ;
    RECT 0.0 188.16 6.24 188.96 ;
    LAYER M3 ;
    RECT 0.0 191.56 6.24 192.36 ;
    LAYER M3 ;
    RECT 0.0 194.96 6.24 195.76 ;
    LAYER M3 ;
    RECT 0.0 198.36 6.24 199.16 ;
    LAYER M3 ;
    RECT 0.0 201.76 6.24 202.56 ;
    LAYER M3 ;
    RECT 0.0 205.16 6.24 205.96 ;
    LAYER M3 ;
    RECT 0.0 208.56 6.24 209.36 ;
    LAYER M3 ;
    RECT 0.0 211.96 6.24 212.76 ;
    LAYER M3 ;
    RECT 0.0 215.36 6.24 216.16 ;
    LAYER M3 ;
    RECT 0.0 218.76 6.24 219.56 ;
    LAYER M3 ;
    RECT 0.0 222.16 6.24 222.96 ;
    LAYER M3 ;
    RECT 0.0 225.56 6.24 226.36 ;
    LAYER M3 ;
    RECT 0.0 228.96 6.24 229.76 ;
    LAYER M3 ;
    RECT 0.0 232.36 6.24 233.16 ;
    LAYER M3 ;
    RECT 0.0 235.76 6.24 236.56 ;
    LAYER M3 ;
    RECT 0.0 239.16 6.24 239.96 ;
    LAYER M3 ;
    RECT 0.0 242.56 6.24 243.36 ;
    LAYER M3 ;
    RECT 0.0 245.96 6.24 246.76 ;
    LAYER M3 ;
    RECT 0.0 249.36 6.24 250.16 ;
    LAYER M3 ;
    RECT 0.0 252.76 6.24 253.56 ;
    LAYER M3 ;
    RECT 0.0 256.16 6.24 256.96 ;
    LAYER M3 ;
    RECT 0.0 259.56 6.24 260.36 ;
    LAYER M3 ;
    RECT 0.0 262.96 6.24 263.76 ;
    LAYER M3 ;
    RECT 0.0 266.36 6.24 267.16 ;
    LAYER M3 ;
    RECT 0.0 269.76 6.24 270.56 ;
    LAYER M3 ;
    RECT 0.0 273.16 6.24 273.96 ;
    LAYER M3 ;
    RECT 0.0 276.56 6.24 277.36 ;
    LAYER M3 ;
    RECT 0.0 279.96 6.24 280.76 ;
    LAYER M3 ;
    RECT 0.0 283.36 6.24 284.16 ;
    LAYER M3 ;
    RECT 0.0 286.76 6.24 287.56 ;
    LAYER M3 ;
    RECT 0.0 290.16 6.24 290.96 ;
    LAYER M3 ;
    RECT 0.0 293.56 6.24 294.36 ;
    LAYER M3 ;
    RECT 0.0 296.96 6.24 297.76 ;
    LAYER M3 ;
    RECT 0.0 300.36 6.24 301.16 ;
    LAYER M3 ;
    RECT 0.0 303.76 6.24 304.56 ;
    LAYER M3 ;
    RECT 0.0 307.16 6.24 307.96 ;
    LAYER M3 ;
    RECT 0.0 310.56 6.24 311.36 ;
    LAYER M3 ;
    RECT 0.0 313.96 6.24 314.76 ;
    LAYER M3 ;
    RECT 0.0 317.36 6.24 318.16 ;
    LAYER M3 ;
    RECT 0.0 320.76 6.24 321.56 ;
    LAYER M3 ;
    RECT 0.0 324.16 6.24 324.96 ;
    LAYER M3 ;
    RECT 0.0 327.56 6.24 328.36 ;
    LAYER M3 ;
    RECT 0.0 330.96 6.24 331.76 ;
    LAYER M3 ;
    RECT 0.0 334.36 6.24 335.16 ;
    LAYER M3 ;
    RECT 0.0 337.76 6.24 338.56 ;
    LAYER M3 ;
    RECT 0.0 341.16 6.24 341.96 ;
    LAYER M3 ;
    RECT 0.0 344.56 6.24 345.36 ;
    LAYER M3 ;
    RECT 0.0 347.96 6.24 348.76 ;
    LAYER M3 ;
    RECT 0.0 351.36 6.24 352.16 ;
    LAYER M3 ;
    RECT 0.0 354.76 6.24 355.56 ;
    LAYER M3 ;
    RECT 0.0 358.16 6.24 358.96 ;
    LAYER M3 ;
    RECT 0.0 361.56 6.24 362.36 ;
    LAYER M3 ;
    RECT 0.0 364.96 6.24 365.76 ;
    LAYER M3 ;
    RECT 0.0 368.36 6.24 369.16 ;
    LAYER M3 ;
    RECT 0.0 371.76 6.24 372.56 ;
    LAYER M3 ;
    RECT 0.0 375.16 6.24 375.96 ;
    LAYER M3 ;
    RECT 0.0 378.56 6.24 379.36 ;
    LAYER M3 ;
    RECT 0.0 381.96 6.24 382.76 ;
    LAYER M3 ;
    RECT 0.0 385.36 6.24 386.16 ;
    LAYER M3 ;
    RECT 0.0 388.76 6.24 389.56 ;
    LAYER M3 ;
    RECT 0.0 392.16 6.24 392.96 ;
    LAYER M3 ;
    RECT 0.0 395.56 6.24 396.36 ;
    LAYER M3 ;
    RECT 0.0 398.96 6.24 399.76 ;
    LAYER M3 ;
    RECT 0.0 402.36 6.24 403.16 ;
    LAYER M3 ;
    RECT 0.0 405.76 6.24 406.56 ;
    LAYER M3 ;
    RECT 0.0 409.16 6.24 409.96 ;
    LAYER M3 ;
    RECT 0.0 412.56 6.24 413.36 ;
    LAYER M3 ;
    RECT 0.0 415.96 6.24 416.76 ;
    LAYER M3 ;
    RECT 0.0 419.36 6.24 420.16 ;
    LAYER M3 ;
    RECT 0.0 422.76 6.24 423.56 ;
    LAYER M3 ;
    RECT 0.0 426.16 6.24 426.96 ;
    LAYER M3 ;
    RECT 0.0 429.56 6.24 430.36 ;
    LAYER M3 ;
    RECT 0.0 432.96 6.24 433.76 ;
    LAYER M3 ;
    RECT 0.0 436.36 6.24 437.16 ;
    LAYER M3 ;
    RECT 0.0 439.76 6.24 440.56 ;
    LAYER M3 ;
    RECT 0.0 443.16 6.24 443.96 ;
    LAYER M3 ;
    RECT 0.0 446.56 6.24 447.36 ;
    LAYER M3 ;
    RECT 0.0 449.96 6.24 450.76 ;
    LAYER M3 ;
    RECT 0.0 453.36 6.24 454.16 ;
    LAYER M3 ;
    RECT 0.0 456.76 6.24 457.56 ;
    LAYER M3 ;
    RECT 0.0 460.16 6.24 460.96 ;
    LAYER M3 ;
    RECT 0.0 463.56 6.24 464.36 ;
    LAYER M3 ;
    RECT 0.0 466.96 6.24 467.76 ;
    LAYER M3 ;
    RECT 0.0 470.36 6.24 471.16 ;
    LAYER M3 ;
    RECT 0.0 473.76 6.24 474.56 ;
    LAYER M3 ;
    RECT 0.0 477.16 6.24 477.96 ;
    LAYER M3 ;
    RECT 0.0 480.56 6.24 481.36 ;
    LAYER M3 ;
    RECT 0.0 483.96 6.24 484.76 ;
    LAYER M3 ;
    RECT 0.0 487.36 6.24 488.16 ;
    LAYER M3 ;
    RECT 0.0 490.76 6.24 491.56 ;
    LAYER M3 ;
    RECT 0.0 494.16 6.24 494.96 ;
    LAYER M3 ;
    RECT 0.0 497.56 6.24 498.36 ;
    LAYER M3 ;
    RECT 0.0 500.96 6.24 501.76 ;
    LAYER M3 ;
    RECT 0.0 504.36 6.24 505.16 ;
    LAYER M3 ;
    RECT 0.0 505.6 6.24 506.0 ;
    LAYER M3 ;
    RECT 0.0 509.0 6.24 509.8 ;
    #gnd fingers
    LAYER M4 ;
    RECT 7.41 510.94 8.21 514.06 ;
    LAYER M4 ;
    RECT 8.61 510.94 9.41 514.06 ;
    LAYER M4 ;
    RECT 12.21 510.94 13.01 514.06 ;
    LAYER M4 ;
    RECT 13.41 510.94 14.21 514.06 ;
    LAYER M4 ;
    RECT 17.01 510.94 17.81 514.06 ;
    LAYER M4 ;
    RECT 18.21 510.94 19.01 514.06 ;
    LAYER M4 ;
    RECT 21.81 510.94 22.61 514.06 ;
    LAYER M4 ;
    RECT 23.01 510.94 23.81 514.06 ;
    LAYER M4 ;
    RECT 26.61 510.94 27.41 514.06 ;
    LAYER M4 ;
    RECT 27.81 510.94 28.61 514.06 ;
    LAYER M4 ;
    RECT 31.41 510.94 32.21 514.06 ;
    LAYER M4 ;
    RECT 32.61 510.94 33.41 514.06 ;
    LAYER M4 ;
    RECT 36.21 510.94 37.01 514.06 ;
    LAYER M4 ;
    RECT 37.41 510.94 38.21 514.06 ;
    LAYER M4 ;
    RECT 41.01 510.94 41.81 514.06 ;
    LAYER M4 ;
    RECT 42.21 510.94 43.01 514.06 ;
    LAYER M4 ;
    RECT 45.81 510.94 46.61 514.06 ;
    LAYER M4 ;
    RECT 47.01 510.94 47.81 514.06 ;
    LAYER M4 ;
    RECT 48.21 510.94 49.01 514.06 ;
    LAYER M4 ;
    RECT 51.81 510.94 52.61 514.06 ;
    LAYER M4 ;
    RECT 53.01 510.94 53.81 514.06 ;
    LAYER M4 ;
    RECT 56.61 510.94 57.41 514.06 ;
    LAYER M4 ;
    RECT 57.81 510.94 58.61 514.06 ;
    LAYER M4 ;
    RECT 61.41 510.94 62.21 514.06 ;
    LAYER M4 ;
    RECT 62.61 510.94 63.41 514.06 ;
    LAYER M4 ;
    RECT 66.21 510.94 67.01 514.06 ;
    LAYER M4 ;
    RECT 67.41 510.94 68.21 514.06 ;
    LAYER M4 ;
    RECT 71.01 510.94 71.81 514.06 ;
    LAYER M4 ;
    RECT 72.21 510.94 73.01 514.06 ;
    LAYER M4 ;
    RECT 75.81 510.94 76.61 514.06 ;
    LAYER M4 ;
    RECT 77.01 510.94 77.81 514.06 ;
    LAYER M4 ;
    RECT 80.61 510.94 81.41 514.06 ;
    LAYER M4 ;
    RECT 81.81 510.94 82.61 514.06 ;
    LAYER M4 ;
    RECT 85.41 510.94 86.21 514.06 ;
    LAYER M4 ;
    RECT 86.61 510.94 87.41 514.06 ;
    LAYER M4 ;
    RECT 89.11 510.94 90.21 514.06 ;
    LAYER M4 ;
    RECT 92.51 510.94 93.61 514.06 ;
    LAYER M4 ;
    RECT 95.91 510.94 97.01 514.06 ;
    LAYER M4 ;
    RECT 99.31 510.94 100.41 514.06 ;
    LAYER M4 ;
    RECT 102.71 510.94 103.81 514.06 ;
    LAYER M4 ;
    RECT 106.11 510.94 107.21 514.06 ;
    LAYER M4 ;
    RECT 109.51 510.94 110.61 514.06 ;
    LAYER M4 ;
    RECT 114.61 510.94 117.41 514.06 ;
    LAYER M4 ;
    RECT 121.41 510.94 124.21 514.06 ;
    LAYER M4 ;
    RECT 128.21 510.94 131.01 514.06 ;
    LAYER M4 ;
    RECT 135.01 510.94 137.81 514.06 ;
    LAYER M4 ;
    RECT 142.25 510.94 143.57 514.06 ;
    LAYER M4 ;
    RECT 146.09 510.94 147.41 514.06 ;
    LAYER M4 ;
    RECT 149.93 510.94 150.39 514.06 ;
    LAYER M4 ;
    RECT 150.79 510.94 151.59 514.06 ;
    LAYER M4 ;
    RECT 153.19 510.94 153.99 514.06 ;
    LAYER M4 ;
    RECT 154.39 510.94 155.19 514.06 ;
    LAYER M4 ;
    RECT 157.99 510.94 158.79 514.06 ;
    LAYER M4 ;
    RECT 159.19 510.94 159.99 514.06 ;
    LAYER M4 ;
    RECT 162.79 510.94 163.59 514.06 ;
    LAYER M4 ;
    RECT 163.99 510.94 164.79 514.06 ;
    LAYER M4 ;
    RECT 167.59 510.94 168.39 514.06 ;
    LAYER M4 ;
    RECT 168.79 510.94 169.59 514.06 ;
    LAYER M4 ;
    RECT 172.39 510.94 173.19 514.06 ;
    LAYER M4 ;
    RECT 173.59 510.94 174.39 514.06 ;
    LAYER M4 ;
    RECT 177.19 510.94 177.99 514.06 ;
    LAYER M4 ;
    RECT 178.39 510.94 179.19 514.06 ;
    LAYER M4 ;
    RECT 181.99 510.94 182.79 514.06 ;
    LAYER M4 ;
    RECT 183.19 510.94 183.99 514.06 ;
    LAYER M4 ;
    RECT 186.79 510.94 187.59 514.06 ;
    LAYER M4 ;
    RECT 187.99 510.94 188.79 514.06 ;
    LAYER M4 ;
    RECT 191.59 510.94 192.39 514.06 ;
    LAYER M4 ;
    RECT 192.79 510.94 193.59 514.06 ;
    LAYER M4 ;
    RECT 193.99 510.94 194.79 514.06 ;
    LAYER M4 ;
    RECT 197.59 510.94 198.39 514.06 ;
    LAYER M4 ;
    RECT 198.79 510.94 199.59 514.06 ;
    LAYER M4 ;
    RECT 202.39 510.94 203.19 514.06 ;
    LAYER M4 ;
    RECT 203.59 510.94 204.39 514.06 ;
    LAYER M4 ;
    RECT 207.19 510.94 207.99 514.06 ;
    LAYER M4 ;
    RECT 208.39 510.94 209.19 514.06 ;
    LAYER M4 ;
    RECT 211.99 510.94 212.79 514.06 ;
    LAYER M4 ;
    RECT 213.19 510.94 213.99 514.06 ;
    LAYER M4 ;
    RECT 216.79 510.94 217.59 514.06 ;
    LAYER M4 ;
    RECT 217.99 510.94 218.79 514.06 ;
    LAYER M4 ;
    RECT 221.59 510.94 222.39 514.06 ;
    LAYER M4 ;
    RECT 222.79 510.94 223.59 514.06 ;
    LAYER M4 ;
    RECT 226.39 510.94 227.19 514.06 ;
    LAYER M4 ;
    RECT 227.59 510.94 228.39 514.06 ;
    LAYER M4 ;
    RECT 231.19 510.94 231.99 514.06 ;
    LAYER M4 ;
    RECT 232.39 510.94 233.19 514.06 ;
    LAYER M4 ;
    RECT 7.41 3.12 9.41 6.24 ;
    LAYER M4 ;
    RECT 12.21 3.12 14.19 6.24 ;
    LAYER M4 ;
    RECT 17.01 3.12 18.41 6.24 ;
    LAYER M4 ;
    RECT 21.81 3.12 23.31 6.24 ;
    LAYER M4 ;
    RECT 27.21 3.12 28.01 6.24 ;
    LAYER M4 ;
    RECT 31.91 3.12 33.41 6.24 ;
    LAYER M4 ;
    RECT 36.21 3.12 38.21 6.24 ;
    LAYER M4 ;
    RECT 41.03 3.12 43.01 6.24 ;
    LAYER M4 ;
    RECT 45.81 3.12 47.21 6.24 ;
    LAYER M4 ;
    RECT 47.61 3.12 49.01 6.24 ;
    LAYER M4 ;
    RECT 51.81 3.12 53.79 6.24 ;
    LAYER M4 ;
    RECT 56.61 3.12 58.61 6.24 ;
    LAYER M4 ;
    RECT 61.41 3.12 62.91 6.24 ;
    LAYER M4 ;
    RECT 66.81 3.12 67.61 6.24 ;
    LAYER M4 ;
    RECT 71.51 3.12 73.01 6.24 ;
    LAYER M4 ;
    RECT 75.81 3.12 77.81 6.24 ;
    LAYER M4 ;
    RECT 80.63 3.12 82.61 6.24 ;
    LAYER M4 ;
    RECT 85.41 3.12 86.71 6.24 ;
    LAYER M4 ;
    RECT 88.81 3.12 89.79 6.24 ;
    LAYER M4 ;
    RECT 94.63 3.12 96.61 6.24 ;
    LAYER M4 ;
    RECT 101.43 3.12 103.39 6.24 ;
    LAYER M4 ;
    RECT 108.23 3.12 110.21 6.24 ;
    LAYER M4 ;
    RECT 115.03 3.12 116.99 6.24 ;
    LAYER M4 ;
    RECT 121.83 3.12 123.81 6.24 ;
    LAYER M4 ;
    RECT 128.63 3.12 130.59 6.24 ;
    LAYER M4 ;
    RECT 135.43 3.12 137.39 6.24 ;
    LAYER M4 ;
    RECT 142.62 3.12 143.57 6.24 ;
    LAYER M4 ;
    RECT 146.09 3.12 147.41 6.24 ;
    LAYER M4 ;
    RECT 150.29 3.12 150.89 6.24 ;
    LAYER M4 ;
    RECT 153.89 3.12 155.19 6.24 ;
    LAYER M4 ;
    RECT 157.99 3.12 159.97 6.24 ;
    LAYER M4 ;
    RECT 162.79 3.12 164.79 6.24 ;
    LAYER M4 ;
    RECT 167.59 3.12 169.09 6.24 ;
    LAYER M4 ;
    RECT 172.99 3.12 173.79 6.24 ;
    LAYER M4 ;
    RECT 177.69 3.12 179.19 6.24 ;
    LAYER M4 ;
    RECT 181.99 3.12 183.99 6.24 ;
    LAYER M4 ;
    RECT 186.81 3.12 188.79 6.24 ;
    LAYER M4 ;
    RECT 191.59 3.12 192.99 6.24 ;
    LAYER M4 ;
    RECT 193.39 3.12 194.79 6.24 ;
    LAYER M4 ;
    RECT 197.59 3.12 199.57 6.24 ;
    LAYER M4 ;
    RECT 202.39 3.12 204.39 6.24 ;
    LAYER M4 ;
    RECT 207.19 3.12 208.69 6.24 ;
    LAYER M4 ;
    RECT 212.59 3.12 213.39 6.24 ;
    LAYER M4 ;
    RECT 217.29 3.12 218.79 6.24 ;
    LAYER M4 ;
    RECT 221.59 3.12 223.59 6.24 ;
    LAYER M4 ;
    RECT 226.41 3.12 228.39 6.24 ;
    LAYER M4 ;
    RECT 231.19 3.12 233.19 6.24 ;
    LAYER M3 ;
    RECT 234.36 12.64 237.48 13.74 ;
    LAYER M3 ;
    RECT 234.36 21.41 237.48 22.21 ;
    LAYER M3 ;
    RECT 234.36 31.13 237.48 32.13 ;
    LAYER M3 ;
    RECT 234.36 32.98 237.48 33.98 ;
    LAYER M3 ;
    RECT 234.36 39.44 237.48 40.44 ;
    LAYER M3 ;
    RECT 234.36 41.29 237.48 42.29 ;
    LAYER M3 ;
    RECT 234.36 54.22 237.48 55.22 ;
    LAYER M3 ;
    RECT 234.36 70.86 237.48 71.66 ;
    LAYER M3 ;
    RECT 234.36 74.26 237.48 75.06 ;
    LAYER M3 ;
    RECT 234.36 77.66 237.48 78.46 ;
    LAYER M3 ;
    RECT 234.36 81.06 237.48 81.86 ;
    LAYER M3 ;
    RECT 234.36 84.46 237.48 85.26 ;
    LAYER M3 ;
    RECT 234.36 87.86 237.48 88.66 ;
    LAYER M3 ;
    RECT 234.36 91.26 237.48 92.06 ;
    LAYER M3 ;
    RECT 234.36 94.66 237.48 95.46 ;
    LAYER M3 ;
    RECT 234.36 98.06 237.48 98.86 ;
    LAYER M3 ;
    RECT 234.36 101.46 237.48 102.26 ;
    LAYER M3 ;
    RECT 234.36 104.86 237.48 105.66 ;
    LAYER M3 ;
    RECT 234.36 108.26 237.48 109.06 ;
    LAYER M3 ;
    RECT 234.36 111.66 237.48 112.46 ;
    LAYER M3 ;
    RECT 234.36 115.06 237.48 115.86 ;
    LAYER M3 ;
    RECT 234.36 118.46 237.48 119.26 ;
    LAYER M3 ;
    RECT 234.36 121.86 237.48 122.66 ;
    LAYER M3 ;
    RECT 234.36 125.26 237.48 126.06 ;
    LAYER M3 ;
    RECT 234.36 128.66 237.48 129.46 ;
    LAYER M3 ;
    RECT 234.36 132.06 237.48 132.86 ;
    LAYER M3 ;
    RECT 234.36 135.46 237.48 136.26 ;
    LAYER M3 ;
    RECT 234.36 138.86 237.48 139.66 ;
    LAYER M3 ;
    RECT 234.36 142.26 237.48 143.06 ;
    LAYER M3 ;
    RECT 234.36 145.66 237.48 146.46 ;
    LAYER M3 ;
    RECT 234.36 149.06 237.48 149.86 ;
    LAYER M3 ;
    RECT 234.36 152.46 237.48 153.26 ;
    LAYER M3 ;
    RECT 234.36 155.86 237.48 156.66 ;
    LAYER M3 ;
    RECT 234.36 159.26 237.48 160.06 ;
    LAYER M3 ;
    RECT 234.36 162.66 237.48 163.46 ;
    LAYER M3 ;
    RECT 234.36 166.06 237.48 166.86 ;
    LAYER M3 ;
    RECT 234.36 169.46 237.48 170.26 ;
    LAYER M3 ;
    RECT 234.36 172.86 237.48 173.66 ;
    LAYER M3 ;
    RECT 234.36 176.26 237.48 177.06 ;
    LAYER M3 ;
    RECT 234.36 179.66 237.48 180.46 ;
    LAYER M3 ;
    RECT 234.36 183.06 237.48 183.86 ;
    LAYER M3 ;
    RECT 234.36 186.46 237.48 187.26 ;
    LAYER M3 ;
    RECT 234.36 189.86 237.48 190.66 ;
    LAYER M3 ;
    RECT 234.36 193.26 237.48 194.06 ;
    LAYER M3 ;
    RECT 234.36 196.66 237.48 197.46 ;
    LAYER M3 ;
    RECT 234.36 200.06 237.48 200.86 ;
    LAYER M3 ;
    RECT 234.36 203.46 237.48 204.26 ;
    LAYER M3 ;
    RECT 234.36 206.86 237.48 207.66 ;
    LAYER M3 ;
    RECT 234.36 210.26 237.48 211.06 ;
    LAYER M3 ;
    RECT 234.36 213.66 237.48 214.46 ;
    LAYER M3 ;
    RECT 234.36 217.06 237.48 217.86 ;
    LAYER M3 ;
    RECT 234.36 220.46 237.48 221.26 ;
    LAYER M3 ;
    RECT 234.36 223.86 237.48 224.66 ;
    LAYER M3 ;
    RECT 234.36 227.26 237.48 228.06 ;
    LAYER M3 ;
    RECT 234.36 230.66 237.48 231.46 ;
    LAYER M3 ;
    RECT 234.36 234.06 237.48 234.86 ;
    LAYER M3 ;
    RECT 234.36 237.46 237.48 238.26 ;
    LAYER M3 ;
    RECT 234.36 240.86 237.48 241.66 ;
    LAYER M3 ;
    RECT 234.36 244.26 237.48 245.06 ;
    LAYER M3 ;
    RECT 234.36 247.66 237.48 248.46 ;
    LAYER M3 ;
    RECT 234.36 251.06 237.48 251.86 ;
    LAYER M3 ;
    RECT 234.36 254.46 237.48 255.26 ;
    LAYER M3 ;
    RECT 234.36 257.86 237.48 258.66 ;
    LAYER M3 ;
    RECT 234.36 261.26 237.48 262.06 ;
    LAYER M3 ;
    RECT 234.36 264.66 237.48 265.46 ;
    LAYER M3 ;
    RECT 234.36 268.06 237.48 268.86 ;
    LAYER M3 ;
    RECT 234.36 271.46 237.48 272.26 ;
    LAYER M3 ;
    RECT 234.36 274.86 237.48 275.66 ;
    LAYER M3 ;
    RECT 234.36 278.26 237.48 279.06 ;
    LAYER M3 ;
    RECT 234.36 281.66 237.48 282.46 ;
    LAYER M3 ;
    RECT 234.36 285.06 237.48 285.86 ;
    LAYER M3 ;
    RECT 234.36 288.46 237.48 289.26 ;
    LAYER M3 ;
    RECT 234.36 291.86 237.48 292.66 ;
    LAYER M3 ;
    RECT 234.36 295.26 237.48 296.06 ;
    LAYER M3 ;
    RECT 234.36 298.66 237.48 299.46 ;
    LAYER M3 ;
    RECT 234.36 302.06 237.48 302.86 ;
    LAYER M3 ;
    RECT 234.36 305.46 237.48 306.26 ;
    LAYER M3 ;
    RECT 234.36 308.86 237.48 309.66 ;
    LAYER M3 ;
    RECT 234.36 312.26 237.48 313.06 ;
    LAYER M3 ;
    RECT 234.36 315.66 237.48 316.46 ;
    LAYER M3 ;
    RECT 234.36 319.06 237.48 319.86 ;
    LAYER M3 ;
    RECT 234.36 322.46 237.48 323.26 ;
    LAYER M3 ;
    RECT 234.36 325.86 237.48 326.66 ;
    LAYER M3 ;
    RECT 234.36 329.26 237.48 330.06 ;
    LAYER M3 ;
    RECT 234.36 332.66 237.48 333.46 ;
    LAYER M3 ;
    RECT 234.36 336.06 237.48 336.86 ;
    LAYER M3 ;
    RECT 234.36 339.46 237.48 340.26 ;
    LAYER M3 ;
    RECT 234.36 342.86 237.48 343.66 ;
    LAYER M3 ;
    RECT 234.36 346.26 237.48 347.06 ;
    LAYER M3 ;
    RECT 234.36 349.66 237.48 350.46 ;
    LAYER M3 ;
    RECT 234.36 353.06 237.48 353.86 ;
    LAYER M3 ;
    RECT 234.36 356.46 237.48 357.26 ;
    LAYER M3 ;
    RECT 234.36 359.86 237.48 360.66 ;
    LAYER M3 ;
    RECT 234.36 363.26 237.48 364.06 ;
    LAYER M3 ;
    RECT 234.36 366.66 237.48 367.46 ;
    LAYER M3 ;
    RECT 234.36 370.06 237.48 370.86 ;
    LAYER M3 ;
    RECT 234.36 373.46 237.48 374.26 ;
    LAYER M3 ;
    RECT 234.36 376.86 237.48 377.66 ;
    LAYER M3 ;
    RECT 234.36 380.26 237.48 381.06 ;
    LAYER M3 ;
    RECT 234.36 383.66 237.48 384.46 ;
    LAYER M3 ;
    RECT 234.36 387.06 237.48 387.86 ;
    LAYER M3 ;
    RECT 234.36 390.46 237.48 391.26 ;
    LAYER M3 ;
    RECT 234.36 393.86 237.48 394.66 ;
    LAYER M3 ;
    RECT 234.36 397.26 237.48 398.06 ;
    LAYER M3 ;
    RECT 234.36 400.66 237.48 401.46 ;
    LAYER M3 ;
    RECT 234.36 404.06 237.48 404.86 ;
    LAYER M3 ;
    RECT 234.36 407.46 237.48 408.26 ;
    LAYER M3 ;
    RECT 234.36 410.86 237.48 411.66 ;
    LAYER M3 ;
    RECT 234.36 414.26 237.48 415.06 ;
    LAYER M3 ;
    RECT 234.36 417.66 237.48 418.46 ;
    LAYER M3 ;
    RECT 234.36 421.06 237.48 421.86 ;
    LAYER M3 ;
    RECT 234.36 424.46 237.48 425.26 ;
    LAYER M3 ;
    RECT 234.36 427.86 237.48 428.66 ;
    LAYER M3 ;
    RECT 234.36 431.26 237.48 432.06 ;
    LAYER M3 ;
    RECT 234.36 434.66 237.48 435.46 ;
    LAYER M3 ;
    RECT 234.36 438.06 237.48 438.86 ;
    LAYER M3 ;
    RECT 234.36 441.46 237.48 442.26 ;
    LAYER M3 ;
    RECT 234.36 444.86 237.48 445.66 ;
    LAYER M3 ;
    RECT 234.36 448.26 237.48 449.06 ;
    LAYER M3 ;
    RECT 234.36 451.66 237.48 452.46 ;
    LAYER M3 ;
    RECT 234.36 455.06 237.48 455.86 ;
    LAYER M3 ;
    RECT 234.36 458.46 237.48 459.26 ;
    LAYER M3 ;
    RECT 234.36 461.86 237.48 462.66 ;
    LAYER M3 ;
    RECT 234.36 465.26 237.48 466.06 ;
    LAYER M3 ;
    RECT 234.36 468.66 237.48 469.46 ;
    LAYER M3 ;
    RECT 234.36 472.06 237.48 472.86 ;
    LAYER M3 ;
    RECT 234.36 475.46 237.48 476.26 ;
    LAYER M3 ;
    RECT 234.36 478.86 237.48 479.66 ;
    LAYER M3 ;
    RECT 234.36 482.26 237.48 483.06 ;
    LAYER M3 ;
    RECT 234.36 485.66 237.48 486.46 ;
    LAYER M3 ;
    RECT 234.36 489.06 237.48 489.86 ;
    LAYER M3 ;
    RECT 234.36 492.46 237.48 493.26 ;
    LAYER M3 ;
    RECT 234.36 495.86 237.48 496.66 ;
    LAYER M3 ;
    RECT 234.36 499.26 237.48 500.06 ;
    LAYER M3 ;
    RECT 234.36 502.66 237.48 503.46 ;
    LAYER M3 ;
    RECT 234.36 506.6 237.48 508.6 ;
    LAYER M3 ;
    RECT 3.12 12.64 6.24 13.74 ;
    LAYER M3 ;
    RECT 3.12 21.41 6.24 22.21 ;
    LAYER M3 ;
    RECT 3.12 31.13 6.24 32.13 ;
    LAYER M3 ;
    RECT 3.12 32.98 6.24 33.98 ;
    LAYER M3 ;
    RECT 3.12 39.44 6.24 40.44 ;
    LAYER M3 ;
    RECT 3.12 41.29 6.24 42.29 ;
    LAYER M3 ;
    RECT 3.12 54.22 6.24 55.22 ;
    LAYER M3 ;
    RECT 3.12 70.86 6.24 71.66 ;
    LAYER M3 ;
    RECT 3.12 74.26 6.24 75.06 ;
    LAYER M3 ;
    RECT 3.12 77.66 6.24 78.46 ;
    LAYER M3 ;
    RECT 3.12 81.06 6.24 81.86 ;
    LAYER M3 ;
    RECT 3.12 84.46 6.24 85.26 ;
    LAYER M3 ;
    RECT 3.12 87.86 6.24 88.66 ;
    LAYER M3 ;
    RECT 3.12 91.26 6.24 92.06 ;
    LAYER M3 ;
    RECT 3.12 94.66 6.24 95.46 ;
    LAYER M3 ;
    RECT 3.12 98.06 6.24 98.86 ;
    LAYER M3 ;
    RECT 3.12 101.46 6.24 102.26 ;
    LAYER M3 ;
    RECT 3.12 104.86 6.24 105.66 ;
    LAYER M3 ;
    RECT 3.12 108.26 6.24 109.06 ;
    LAYER M3 ;
    RECT 3.12 111.66 6.24 112.46 ;
    LAYER M3 ;
    RECT 3.12 115.06 6.24 115.86 ;
    LAYER M3 ;
    RECT 3.12 118.46 6.24 119.26 ;
    LAYER M3 ;
    RECT 3.12 121.86 6.24 122.66 ;
    LAYER M3 ;
    RECT 3.12 125.26 6.24 126.06 ;
    LAYER M3 ;
    RECT 3.12 128.66 6.24 129.46 ;
    LAYER M3 ;
    RECT 3.12 132.06 6.24 132.86 ;
    LAYER M3 ;
    RECT 3.12 135.46 6.24 136.26 ;
    LAYER M3 ;
    RECT 3.12 138.86 6.24 139.66 ;
    LAYER M3 ;
    RECT 3.12 142.26 6.24 143.06 ;
    LAYER M3 ;
    RECT 3.12 145.66 6.24 146.46 ;
    LAYER M3 ;
    RECT 3.12 149.06 6.24 149.86 ;
    LAYER M3 ;
    RECT 3.12 152.46 6.24 153.26 ;
    LAYER M3 ;
    RECT 3.12 155.86 6.24 156.66 ;
    LAYER M3 ;
    RECT 3.12 159.26 6.24 160.06 ;
    LAYER M3 ;
    RECT 3.12 162.66 6.24 163.46 ;
    LAYER M3 ;
    RECT 3.12 166.06 6.24 166.86 ;
    LAYER M3 ;
    RECT 3.12 169.46 6.24 170.26 ;
    LAYER M3 ;
    RECT 3.12 172.86 6.24 173.66 ;
    LAYER M3 ;
    RECT 3.12 176.26 6.24 177.06 ;
    LAYER M3 ;
    RECT 3.12 179.66 6.24 180.46 ;
    LAYER M3 ;
    RECT 3.12 183.06 6.24 183.86 ;
    LAYER M3 ;
    RECT 3.12 186.46 6.24 187.26 ;
    LAYER M3 ;
    RECT 3.12 189.86 6.24 190.66 ;
    LAYER M3 ;
    RECT 3.12 193.26 6.24 194.06 ;
    LAYER M3 ;
    RECT 3.12 196.66 6.24 197.46 ;
    LAYER M3 ;
    RECT 3.12 200.06 6.24 200.86 ;
    LAYER M3 ;
    RECT 3.12 203.46 6.24 204.26 ;
    LAYER M3 ;
    RECT 3.12 206.86 6.24 207.66 ;
    LAYER M3 ;
    RECT 3.12 210.26 6.24 211.06 ;
    LAYER M3 ;
    RECT 3.12 213.66 6.24 214.46 ;
    LAYER M3 ;
    RECT 3.12 217.06 6.24 217.86 ;
    LAYER M3 ;
    RECT 3.12 220.46 6.24 221.26 ;
    LAYER M3 ;
    RECT 3.12 223.86 6.24 224.66 ;
    LAYER M3 ;
    RECT 3.12 227.26 6.24 228.06 ;
    LAYER M3 ;
    RECT 3.12 230.66 6.24 231.46 ;
    LAYER M3 ;
    RECT 3.12 234.06 6.24 234.86 ;
    LAYER M3 ;
    RECT 3.12 237.46 6.24 238.26 ;
    LAYER M3 ;
    RECT 3.12 240.86 6.24 241.66 ;
    LAYER M3 ;
    RECT 3.12 244.26 6.24 245.06 ;
    LAYER M3 ;
    RECT 3.12 247.66 6.24 248.46 ;
    LAYER M3 ;
    RECT 3.12 251.06 6.24 251.86 ;
    LAYER M3 ;
    RECT 3.12 254.46 6.24 255.26 ;
    LAYER M3 ;
    RECT 3.12 257.86 6.24 258.66 ;
    LAYER M3 ;
    RECT 3.12 261.26 6.24 262.06 ;
    LAYER M3 ;
    RECT 3.12 264.66 6.24 265.46 ;
    LAYER M3 ;
    RECT 3.12 268.06 6.24 268.86 ;
    LAYER M3 ;
    RECT 3.12 271.46 6.24 272.26 ;
    LAYER M3 ;
    RECT 3.12 274.86 6.24 275.66 ;
    LAYER M3 ;
    RECT 3.12 278.26 6.24 279.06 ;
    LAYER M3 ;
    RECT 3.12 281.66 6.24 282.46 ;
    LAYER M3 ;
    RECT 3.12 285.06 6.24 285.86 ;
    LAYER M3 ;
    RECT 3.12 288.46 6.24 289.26 ;
    LAYER M3 ;
    RECT 3.12 291.86 6.24 292.66 ;
    LAYER M3 ;
    RECT 3.12 295.26 6.24 296.06 ;
    LAYER M3 ;
    RECT 3.12 298.66 6.24 299.46 ;
    LAYER M3 ;
    RECT 3.12 302.06 6.24 302.86 ;
    LAYER M3 ;
    RECT 3.12 305.46 6.24 306.26 ;
    LAYER M3 ;
    RECT 3.12 308.86 6.24 309.66 ;
    LAYER M3 ;
    RECT 3.12 312.26 6.24 313.06 ;
    LAYER M3 ;
    RECT 3.12 315.66 6.24 316.46 ;
    LAYER M3 ;
    RECT 3.12 319.06 6.24 319.86 ;
    LAYER M3 ;
    RECT 3.12 322.46 6.24 323.26 ;
    LAYER M3 ;
    RECT 3.12 325.86 6.24 326.66 ;
    LAYER M3 ;
    RECT 3.12 329.26 6.24 330.06 ;
    LAYER M3 ;
    RECT 3.12 332.66 6.24 333.46 ;
    LAYER M3 ;
    RECT 3.12 336.06 6.24 336.86 ;
    LAYER M3 ;
    RECT 3.12 339.46 6.24 340.26 ;
    LAYER M3 ;
    RECT 3.12 342.86 6.24 343.66 ;
    LAYER M3 ;
    RECT 3.12 346.26 6.24 347.06 ;
    LAYER M3 ;
    RECT 3.12 349.66 6.24 350.46 ;
    LAYER M3 ;
    RECT 3.12 353.06 6.24 353.86 ;
    LAYER M3 ;
    RECT 3.12 356.46 6.24 357.26 ;
    LAYER M3 ;
    RECT 3.12 359.86 6.24 360.66 ;
    LAYER M3 ;
    RECT 3.12 363.26 6.24 364.06 ;
    LAYER M3 ;
    RECT 3.12 366.66 6.24 367.46 ;
    LAYER M3 ;
    RECT 3.12 370.06 6.24 370.86 ;
    LAYER M3 ;
    RECT 3.12 373.46 6.24 374.26 ;
    LAYER M3 ;
    RECT 3.12 376.86 6.24 377.66 ;
    LAYER M3 ;
    RECT 3.12 380.26 6.24 381.06 ;
    LAYER M3 ;
    RECT 3.12 383.66 6.24 384.46 ;
    LAYER M3 ;
    RECT 3.12 387.06 6.24 387.86 ;
    LAYER M3 ;
    RECT 3.12 390.46 6.24 391.26 ;
    LAYER M3 ;
    RECT 3.12 393.86 6.24 394.66 ;
    LAYER M3 ;
    RECT 3.12 397.26 6.24 398.06 ;
    LAYER M3 ;
    RECT 3.12 400.66 6.24 401.46 ;
    LAYER M3 ;
    RECT 3.12 404.06 6.24 404.86 ;
    LAYER M3 ;
    RECT 3.12 407.46 6.24 408.26 ;
    LAYER M3 ;
    RECT 3.12 410.86 6.24 411.66 ;
    LAYER M3 ;
    RECT 3.12 414.26 6.24 415.06 ;
    LAYER M3 ;
    RECT 3.12 417.66 6.24 418.46 ;
    LAYER M3 ;
    RECT 3.12 421.06 6.24 421.86 ;
    LAYER M3 ;
    RECT 3.12 424.46 6.24 425.26 ;
    LAYER M3 ;
    RECT 3.12 427.86 6.24 428.66 ;
    LAYER M3 ;
    RECT 3.12 431.26 6.24 432.06 ;
    LAYER M3 ;
    RECT 3.12 434.66 6.24 435.46 ;
    LAYER M3 ;
    RECT 3.12 438.06 6.24 438.86 ;
    LAYER M3 ;
    RECT 3.12 441.46 6.24 442.26 ;
    LAYER M3 ;
    RECT 3.12 444.86 6.24 445.66 ;
    LAYER M3 ;
    RECT 3.12 448.26 6.24 449.06 ;
    LAYER M3 ;
    RECT 3.12 451.66 6.24 452.46 ;
    LAYER M3 ;
    RECT 3.12 455.06 6.24 455.86 ;
    LAYER M3 ;
    RECT 3.12 458.46 6.24 459.26 ;
    LAYER M3 ;
    RECT 3.12 461.86 6.24 462.66 ;
    LAYER M3 ;
    RECT 3.12 465.26 6.24 466.06 ;
    LAYER M3 ;
    RECT 3.12 468.66 6.24 469.46 ;
    LAYER M3 ;
    RECT 3.12 472.06 6.24 472.86 ;
    LAYER M3 ;
    RECT 3.12 475.46 6.24 476.26 ;
    LAYER M3 ;
    RECT 3.12 478.86 6.24 479.66 ;
    LAYER M3 ;
    RECT 3.12 482.26 6.24 483.06 ;
    LAYER M3 ;
    RECT 3.12 485.66 6.24 486.46 ;
    LAYER M3 ;
    RECT 3.12 489.06 6.24 489.86 ;
    LAYER M3 ;
    RECT 3.12 492.46 6.24 493.26 ;
    LAYER M3 ;
    RECT 3.12 495.86 6.24 496.66 ;
    LAYER M3 ;
    RECT 3.12 499.26 6.24 500.06 ;
    LAYER M3 ;
    RECT 3.12 502.66 6.24 503.46 ;
    LAYER M3 ;
    RECT 3.12 506.6 6.24 508.6 ;
    #ring waffles
    LAYER V3 ;
    RECT 3.12 512.06 5.12 514.06 ;
    LAYER V3 ;
    RECT 235.48 512.06 237.48 514.06 ;
    LAYER V3 ;
    RECT 3.12 3.12 5.12 5.12 ;
    LAYER V3 ;
    RECT 235.48 3.12 237.48 5.12 ;
    LAYER V3 ;
    RECT 0.0 515.18 2.0 517.18 ;
    LAYER V3 ;
    RECT 238.6 515.18 240.6 517.18 ;
    LAYER V3 ;
    RECT 0.0 0.0 2.0 2.0 ;
    LAYER V3 ;
    RECT 238.6 0.0 240.6 2.0 ;
    #finger waffles
    LAYER V3 ;
    RECT 7.41 512.06 8.21 514.06 ;
    LAYER V3 ;
    RECT 8.61 512.06 9.41 514.06 ;
    LAYER V3 ;
    RECT 9.81 515.18 11.81 517.18 ;
    LAYER V3 ;
    RECT 12.21 512.06 13.01 514.06 ;
    LAYER V3 ;
    RECT 13.41 512.06 14.21 514.06 ;
    LAYER V3 ;
    RECT 14.61 515.18 16.61 517.18 ;
    LAYER V3 ;
    RECT 17.01 512.06 17.81 514.06 ;
    LAYER V3 ;
    RECT 18.21 512.06 19.01 514.06 ;
    LAYER V3 ;
    RECT 19.41 515.18 21.41 517.18 ;
    LAYER V3 ;
    RECT 21.81 512.06 22.61 514.06 ;
    LAYER V3 ;
    RECT 23.01 512.06 23.81 514.06 ;
    LAYER V3 ;
    RECT 24.21 515.18 26.21 517.18 ;
    LAYER V3 ;
    RECT 26.61 512.06 27.41 514.06 ;
    LAYER V3 ;
    RECT 27.81 512.06 28.61 514.06 ;
    LAYER V3 ;
    RECT 29.01 515.18 31.01 517.18 ;
    LAYER V3 ;
    RECT 31.41 512.06 32.21 514.06 ;
    LAYER V3 ;
    RECT 32.61 512.06 33.41 514.06 ;
    LAYER V3 ;
    RECT 33.81 515.18 35.81 517.18 ;
    LAYER V3 ;
    RECT 36.21 512.06 37.01 514.06 ;
    LAYER V3 ;
    RECT 37.41 512.06 38.21 514.06 ;
    LAYER V3 ;
    RECT 38.61 515.18 40.61 517.18 ;
    LAYER V3 ;
    RECT 41.01 512.06 41.81 514.06 ;
    LAYER V3 ;
    RECT 42.21 512.06 43.01 514.06 ;
    LAYER V3 ;
    RECT 43.41 515.18 45.41 517.18 ;
    LAYER V3 ;
    RECT 45.81 512.06 46.61 514.06 ;
    LAYER V3 ;
    RECT 47.01 512.06 47.81 514.06 ;
    LAYER V3 ;
    RECT 48.21 512.06 49.01 514.06 ;
    LAYER V3 ;
    RECT 49.41 515.18 51.41 517.18 ;
    LAYER V3 ;
    RECT 51.81 512.06 52.61 514.06 ;
    LAYER V3 ;
    RECT 53.01 512.06 53.81 514.06 ;
    LAYER V3 ;
    RECT 54.21 515.18 56.21 517.18 ;
    LAYER V3 ;
    RECT 56.61 512.06 57.41 514.06 ;
    LAYER V3 ;
    RECT 57.81 512.06 58.61 514.06 ;
    LAYER V3 ;
    RECT 59.01 515.18 61.01 517.18 ;
    LAYER V3 ;
    RECT 61.41 512.06 62.21 514.06 ;
    LAYER V3 ;
    RECT 62.61 512.06 63.41 514.06 ;
    LAYER V3 ;
    RECT 63.81 515.18 65.81 517.18 ;
    LAYER V3 ;
    RECT 66.21 512.06 67.01 514.06 ;
    LAYER V3 ;
    RECT 67.41 512.06 68.21 514.06 ;
    LAYER V3 ;
    RECT 68.61 515.18 70.61 517.18 ;
    LAYER V3 ;
    RECT 71.01 512.06 71.81 514.06 ;
    LAYER V3 ;
    RECT 72.21 512.06 73.01 514.06 ;
    LAYER V3 ;
    RECT 73.41 515.18 75.41 517.18 ;
    LAYER V3 ;
    RECT 75.81 512.06 76.61 514.06 ;
    LAYER V3 ;
    RECT 77.01 512.06 77.81 514.06 ;
    LAYER V3 ;
    RECT 78.21 515.18 80.21 517.18 ;
    LAYER V3 ;
    RECT 80.61 512.06 81.41 514.06 ;
    LAYER V3 ;
    RECT 81.81 512.06 82.61 514.06 ;
    LAYER V3 ;
    RECT 83.01 515.18 85.01 517.18 ;
    LAYER V3 ;
    RECT 85.41 512.06 86.21 514.06 ;
    LAYER V3 ;
    RECT 86.61 512.06 87.41 514.06 ;
    LAYER V3 ;
    RECT 87.81 515.18 88.61 517.18 ;
    LAYER V3 ;
    RECT 89.11 512.06 90.21 514.06 ;
    LAYER V3 ;
    RECT 90.81 515.18 91.91 517.18 ;
    LAYER V3 ;
    RECT 92.51 512.06 93.61 514.06 ;
    LAYER V3 ;
    RECT 94.21 515.18 95.31 517.18 ;
    LAYER V3 ;
    RECT 95.91 512.06 97.01 514.06 ;
    LAYER V3 ;
    RECT 97.61 515.18 98.71 517.18 ;
    LAYER V3 ;
    RECT 99.31 512.06 100.41 514.06 ;
    LAYER V3 ;
    RECT 101.01 515.18 102.11 517.18 ;
    LAYER V3 ;
    RECT 102.71 512.06 103.81 514.06 ;
    LAYER V3 ;
    RECT 104.41 515.18 105.51 517.18 ;
    LAYER V3 ;
    RECT 106.11 512.06 107.21 514.06 ;
    LAYER V3 ;
    RECT 107.81 515.18 108.91 517.18 ;
    LAYER V3 ;
    RECT 109.51 512.06 110.61 514.06 ;
    LAYER V3 ;
    RECT 111.21 515.18 114.01 517.18 ;
    LAYER V3 ;
    RECT 114.61 512.06 117.41 514.06 ;
    LAYER V3 ;
    RECT 118.01 515.18 120.81 517.18 ;
    LAYER V3 ;
    RECT 121.41 512.06 124.21 514.06 ;
    LAYER V3 ;
    RECT 124.81 515.18 127.61 517.18 ;
    LAYER V3 ;
    RECT 128.21 512.06 131.01 514.06 ;
    LAYER V3 ;
    RECT 131.61 515.18 134.41 517.18 ;
    LAYER V3 ;
    RECT 135.01 512.06 137.81 514.06 ;
    LAYER V3 ;
    RECT 138.41 515.18 141.65 517.18 ;
    LAYER V3 ;
    RECT 142.25 512.06 143.57 514.06 ;
    LAYER V3 ;
    RECT 144.17 515.18 145.49 517.18 ;
    LAYER V3 ;
    RECT 146.09 512.06 147.41 514.06 ;
    LAYER V3 ;
    RECT 148.01 515.18 149.33 517.18 ;
    LAYER V3 ;
    RECT 149.93 512.06 150.39 514.06 ;
    LAYER V3 ;
    RECT 150.79 512.06 151.59 514.06 ;
    LAYER V3 ;
    RECT 151.99 515.18 152.79 517.18 ;
    LAYER V3 ;
    RECT 153.19 512.06 153.99 514.06 ;
    LAYER V3 ;
    RECT 154.39 512.06 155.19 514.06 ;
    LAYER V3 ;
    RECT 155.59 515.18 157.59 517.18 ;
    LAYER V3 ;
    RECT 157.99 512.06 158.79 514.06 ;
    LAYER V3 ;
    RECT 159.19 512.06 159.99 514.06 ;
    LAYER V3 ;
    RECT 160.39 515.18 162.39 517.18 ;
    LAYER V3 ;
    RECT 162.79 512.06 163.59 514.06 ;
    LAYER V3 ;
    RECT 163.99 512.06 164.79 514.06 ;
    LAYER V3 ;
    RECT 165.19 515.18 167.19 517.18 ;
    LAYER V3 ;
    RECT 167.59 512.06 168.39 514.06 ;
    LAYER V3 ;
    RECT 168.79 512.06 169.59 514.06 ;
    LAYER V3 ;
    RECT 169.99 515.18 171.99 517.18 ;
    LAYER V3 ;
    RECT 172.39 512.06 173.19 514.06 ;
    LAYER V3 ;
    RECT 173.59 512.06 174.39 514.06 ;
    LAYER V3 ;
    RECT 174.79 515.18 176.79 517.18 ;
    LAYER V3 ;
    RECT 177.19 512.06 177.99 514.06 ;
    LAYER V3 ;
    RECT 178.39 512.06 179.19 514.06 ;
    LAYER V3 ;
    RECT 179.59 515.18 181.59 517.18 ;
    LAYER V3 ;
    RECT 181.99 512.06 182.79 514.06 ;
    LAYER V3 ;
    RECT 183.19 512.06 183.99 514.06 ;
    LAYER V3 ;
    RECT 184.39 515.18 186.39 517.18 ;
    LAYER V3 ;
    RECT 186.79 512.06 187.59 514.06 ;
    LAYER V3 ;
    RECT 187.99 512.06 188.79 514.06 ;
    LAYER V3 ;
    RECT 189.19 515.18 191.19 517.18 ;
    LAYER V3 ;
    RECT 191.59 512.06 192.39 514.06 ;
    LAYER V3 ;
    RECT 192.79 512.06 193.59 514.06 ;
    LAYER V3 ;
    RECT 193.99 512.06 194.79 514.06 ;
    LAYER V3 ;
    RECT 195.19 515.18 197.19 517.18 ;
    LAYER V3 ;
    RECT 197.59 512.06 198.39 514.06 ;
    LAYER V3 ;
    RECT 198.79 512.06 199.59 514.06 ;
    LAYER V3 ;
    RECT 199.99 515.18 201.99 517.18 ;
    LAYER V3 ;
    RECT 202.39 512.06 203.19 514.06 ;
    LAYER V3 ;
    RECT 203.59 512.06 204.39 514.06 ;
    LAYER V3 ;
    RECT 204.79 515.18 206.79 517.18 ;
    LAYER V3 ;
    RECT 207.19 512.06 207.99 514.06 ;
    LAYER V3 ;
    RECT 208.39 512.06 209.19 514.06 ;
    LAYER V3 ;
    RECT 209.59 515.18 211.59 517.18 ;
    LAYER V3 ;
    RECT 211.99 512.06 212.79 514.06 ;
    LAYER V3 ;
    RECT 213.19 512.06 213.99 514.06 ;
    LAYER V3 ;
    RECT 214.39 515.18 216.39 517.18 ;
    LAYER V3 ;
    RECT 216.79 512.06 217.59 514.06 ;
    LAYER V3 ;
    RECT 217.99 512.06 218.79 514.06 ;
    LAYER V3 ;
    RECT 219.19 515.18 221.19 517.18 ;
    LAYER V3 ;
    RECT 221.59 512.06 222.39 514.06 ;
    LAYER V3 ;
    RECT 222.79 512.06 223.59 514.06 ;
    LAYER V3 ;
    RECT 223.99 515.18 225.99 517.18 ;
    LAYER V3 ;
    RECT 226.39 512.06 227.19 514.06 ;
    LAYER V3 ;
    RECT 227.59 512.06 228.39 514.06 ;
    LAYER V3 ;
    RECT 228.79 515.18 230.79 517.18 ;
    LAYER V3 ;
    RECT 231.19 512.06 231.99 514.06 ;
    LAYER V3 ;
    RECT 232.39 512.06 233.19 514.06 ;
    LAYER V3 ;
    RECT 7.41 3.12 9.41 5.12 ;
    LAYER V3 ;
    RECT 9.81 0.0 11.79 2.0 ;
    LAYER V3 ;
    RECT 12.21 3.12 14.19 5.12 ;
    LAYER V3 ;
    RECT 14.61 0.0 16.59 2.0 ;
    LAYER V3 ;
    RECT 17.01 3.12 18.41 5.12 ;
    LAYER V3 ;
    RECT 19.81 0.0 21.41 2.0 ;
    LAYER V3 ;
    RECT 21.81 3.12 23.31 5.12 ;
    LAYER V3 ;
    RECT 24.71 0.0 25.71 2.0 ;
    LAYER V3 ;
    RECT 27.21 3.12 28.01 5.12 ;
    LAYER V3 ;
    RECT 29.51 0.0 30.51 2.0 ;
    LAYER V3 ;
    RECT 31.91 3.12 33.41 5.12 ;
    LAYER V3 ;
    RECT 33.84 0.0 35.81 2.0 ;
    LAYER V3 ;
    RECT 36.21 3.12 38.21 5.12 ;
    LAYER V3 ;
    RECT 38.63 0.0 40.61 2.0 ;
    LAYER V3 ;
    RECT 41.03 3.12 43.01 5.12 ;
    LAYER V3 ;
    RECT 43.43 0.0 45.41 2.0 ;
    LAYER V3 ;
    RECT 45.81 3.12 47.21 5.12 ;
    LAYER V3 ;
    RECT 47.61 3.12 49.01 5.12 ;
    LAYER V3 ;
    RECT 49.41 0.0 51.39 2.0 ;
    LAYER V3 ;
    RECT 51.81 3.12 53.79 5.12 ;
    LAYER V3 ;
    RECT 54.21 0.0 56.19 2.0 ;
    LAYER V3 ;
    RECT 56.61 3.12 58.61 5.12 ;
    LAYER V3 ;
    RECT 59.01 0.0 60.98 2.0 ;
    LAYER V3 ;
    RECT 61.41 3.12 62.91 5.12 ;
    LAYER V3 ;
    RECT 64.31 0.0 65.31 2.0 ;
    LAYER V3 ;
    RECT 66.81 3.12 67.61 5.12 ;
    LAYER V3 ;
    RECT 69.11 0.0 70.11 2.0 ;
    LAYER V3 ;
    RECT 71.51 3.12 73.01 5.12 ;
    LAYER V3 ;
    RECT 73.44 0.0 75.41 2.0 ;
    LAYER V3 ;
    RECT 75.81 3.12 77.81 5.12 ;
    LAYER V3 ;
    RECT 78.23 0.0 80.21 2.0 ;
    LAYER V3 ;
    RECT 80.63 3.12 82.61 5.12 ;
    LAYER V3 ;
    RECT 83.03 0.0 85.01 2.0 ;
    LAYER V3 ;
    RECT 85.41 3.12 86.71 5.12 ;
    LAYER V3 ;
    RECT 87.21 0.0 88.01 2.0 ;
    LAYER V3 ;
    RECT 88.81 3.12 89.79 5.12 ;
    LAYER V3 ;
    RECT 91.23 0.0 93.19 2.0 ;
    LAYER V3 ;
    RECT 94.63 3.12 96.61 5.12 ;
    LAYER V3 ;
    RECT 98.01 0.0 99.99 2.0 ;
    LAYER V3 ;
    RECT 101.43 3.12 103.39 5.12 ;
    LAYER V3 ;
    RECT 104.83 0.0 106.79 2.0 ;
    LAYER V3 ;
    RECT 108.23 3.12 110.21 5.12 ;
    LAYER V3 ;
    RECT 111.61 0.0 113.59 2.0 ;
    LAYER V3 ;
    RECT 115.03 3.12 116.99 5.12 ;
    LAYER V3 ;
    RECT 118.43 0.0 120.39 2.0 ;
    LAYER V3 ;
    RECT 121.83 3.12 123.81 5.12 ;
    LAYER V3 ;
    RECT 125.21 0.0 127.19 2.0 ;
    LAYER V3 ;
    RECT 128.63 3.12 130.59 5.12 ;
    LAYER V3 ;
    RECT 132.03 0.0 133.99 2.0 ;
    LAYER V3 ;
    RECT 135.43 3.12 137.39 5.12 ;
    LAYER V3 ;
    RECT 138.83 0.0 140.83 2.0 ;
    LAYER V3 ;
    RECT 142.62 3.12 143.57 5.12 ;
    LAYER V3 ;
    RECT 145.01 0.0 145.61 2.0 ;
    LAYER V3 ;
    RECT 146.09 3.12 147.41 5.12 ;
    LAYER V3 ;
    RECT 148.01 0.0 148.87 2.0 ;
    LAYER V3 ;
    RECT 150.29 3.12 150.89 5.12 ;
    LAYER V3 ;
    RECT 153.89 3.12 155.19 5.12 ;
    LAYER V3 ;
    RECT 155.59 0.0 157.57 2.0 ;
    LAYER V3 ;
    RECT 157.99 3.12 159.97 5.12 ;
    LAYER V3 ;
    RECT 160.39 0.0 162.37 2.0 ;
    LAYER V3 ;
    RECT 162.79 3.12 164.79 5.12 ;
    LAYER V3 ;
    RECT 165.19 0.0 167.16 2.0 ;
    LAYER V3 ;
    RECT 167.59 3.12 169.09 5.12 ;
    LAYER V3 ;
    RECT 170.49 0.0 171.49 2.0 ;
    LAYER V3 ;
    RECT 172.99 3.12 173.79 5.12 ;
    LAYER V3 ;
    RECT 175.29 0.0 176.29 2.0 ;
    LAYER V3 ;
    RECT 177.69 3.12 179.19 5.12 ;
    LAYER V3 ;
    RECT 179.62 0.0 181.59 2.0 ;
    LAYER V3 ;
    RECT 181.99 3.12 183.99 5.12 ;
    LAYER V3 ;
    RECT 184.41 0.0 186.39 2.0 ;
    LAYER V3 ;
    RECT 186.81 3.12 188.79 5.12 ;
    LAYER V3 ;
    RECT 189.21 0.0 191.19 2.0 ;
    LAYER V3 ;
    RECT 191.59 3.12 192.99 5.12 ;
    LAYER V3 ;
    RECT 193.39 3.12 194.79 5.12 ;
    LAYER V3 ;
    RECT 195.19 0.0 197.17 2.0 ;
    LAYER V3 ;
    RECT 197.59 3.12 199.57 5.12 ;
    LAYER V3 ;
    RECT 199.99 0.0 201.97 2.0 ;
    LAYER V3 ;
    RECT 202.39 3.12 204.39 5.12 ;
    LAYER V3 ;
    RECT 204.79 0.0 206.76 2.0 ;
    LAYER V3 ;
    RECT 207.19 3.12 208.69 5.12 ;
    LAYER V3 ;
    RECT 210.09 0.0 211.09 2.0 ;
    LAYER V3 ;
    RECT 212.59 3.12 213.39 5.12 ;
    LAYER V3 ;
    RECT 214.89 0.0 215.89 2.0 ;
    LAYER V3 ;
    RECT 217.29 3.12 218.79 5.12 ;
    LAYER V3 ;
    RECT 219.21 0.0 221.19 2.0 ;
    LAYER V3 ;
    RECT 221.59 3.12 223.59 5.12 ;
    LAYER V3 ;
    RECT 224.01 0.0 225.99 2.0 ;
    LAYER V3 ;
    RECT 226.41 3.12 228.39 5.12 ;
    LAYER V3 ;
    RECT 228.81 0.0 230.79 2.0 ;
    LAYER V3 ;
    RECT 231.19 3.12 233.19 5.12 ;
    LAYER V3 ;
    RECT 238.6 7.94 240.6 9.14 ;
    LAYER V3 ;
    RECT 235.48 12.64 237.48 13.74 ;
    LAYER V3 ;
    RECT 238.6 17.26 240.6 18.46 ;
    LAYER V3 ;
    RECT 235.48 21.41 237.48 22.21 ;
    LAYER V3 ;
    RECT 238.6 25.81 240.6 27.81 ;
    LAYER V3 ;
    RECT 235.48 31.13 237.48 32.13 ;
    LAYER V3 ;
    RECT 235.48 32.98 237.48 33.98 ;
    LAYER V3 ;
    RECT 238.6 35.91 240.6 36.91 ;
    LAYER V3 ;
    RECT 235.48 39.44 237.48 40.44 ;
    LAYER V3 ;
    RECT 235.48 41.29 237.48 42.29 ;
    LAYER V3 ;
    RECT 238.6 50.24 240.6 51.24 ;
    LAYER V3 ;
    RECT 235.48 54.22 237.48 55.22 ;
    LAYER V3 ;
    RECT 238.6 57.02 240.6 58.02 ;
    LAYER V3 ;
    RECT 238.6 60.6 240.6 61.6 ;
    LAYER V3 ;
    RECT 238.6 62.45 240.6 63.45 ;
    LAYER V3 ;
    RECT 238.6 69.16 240.6 69.96 ;
    LAYER V3 ;
    RECT 235.48 70.86 237.48 71.66 ;
    LAYER V3 ;
    RECT 238.6 72.56 240.6 73.36 ;
    LAYER V3 ;
    RECT 235.48 74.26 237.48 75.06 ;
    LAYER V3 ;
    RECT 238.6 75.96 240.6 76.76 ;
    LAYER V3 ;
    RECT 235.48 77.66 237.48 78.46 ;
    LAYER V3 ;
    RECT 238.6 79.36 240.6 80.16 ;
    LAYER V3 ;
    RECT 235.48 81.06 237.48 81.86 ;
    LAYER V3 ;
    RECT 238.6 82.76 240.6 83.56 ;
    LAYER V3 ;
    RECT 235.48 84.46 237.48 85.26 ;
    LAYER V3 ;
    RECT 238.6 86.16 240.6 86.96 ;
    LAYER V3 ;
    RECT 235.48 87.86 237.48 88.66 ;
    LAYER V3 ;
    RECT 238.6 89.56 240.6 90.36 ;
    LAYER V3 ;
    RECT 235.48 91.26 237.48 92.06 ;
    LAYER V3 ;
    RECT 238.6 92.96 240.6 93.76 ;
    LAYER V3 ;
    RECT 235.48 94.66 237.48 95.46 ;
    LAYER V3 ;
    RECT 238.6 96.36 240.6 97.16 ;
    LAYER V3 ;
    RECT 235.48 98.06 237.48 98.86 ;
    LAYER V3 ;
    RECT 238.6 99.76 240.6 100.56 ;
    LAYER V3 ;
    RECT 235.48 101.46 237.48 102.26 ;
    LAYER V3 ;
    RECT 238.6 103.16 240.6 103.96 ;
    LAYER V3 ;
    RECT 235.48 104.86 237.48 105.66 ;
    LAYER V3 ;
    RECT 238.6 106.56 240.6 107.36 ;
    LAYER V3 ;
    RECT 235.48 108.26 237.48 109.06 ;
    LAYER V3 ;
    RECT 238.6 109.96 240.6 110.76 ;
    LAYER V3 ;
    RECT 235.48 111.66 237.48 112.46 ;
    LAYER V3 ;
    RECT 238.6 113.36 240.6 114.16 ;
    LAYER V3 ;
    RECT 235.48 115.06 237.48 115.86 ;
    LAYER V3 ;
    RECT 238.6 116.76 240.6 117.56 ;
    LAYER V3 ;
    RECT 235.48 118.46 237.48 119.26 ;
    LAYER V3 ;
    RECT 238.6 120.16 240.6 120.96 ;
    LAYER V3 ;
    RECT 235.48 121.86 237.48 122.66 ;
    LAYER V3 ;
    RECT 238.6 123.56 240.6 124.36 ;
    LAYER V3 ;
    RECT 235.48 125.26 237.48 126.06 ;
    LAYER V3 ;
    RECT 238.6 126.96 240.6 127.76 ;
    LAYER V3 ;
    RECT 235.48 128.66 237.48 129.46 ;
    LAYER V3 ;
    RECT 238.6 130.36 240.6 131.16 ;
    LAYER V3 ;
    RECT 235.48 132.06 237.48 132.86 ;
    LAYER V3 ;
    RECT 238.6 133.76 240.6 134.56 ;
    LAYER V3 ;
    RECT 235.48 135.46 237.48 136.26 ;
    LAYER V3 ;
    RECT 238.6 137.16 240.6 137.96 ;
    LAYER V3 ;
    RECT 235.48 138.86 237.48 139.66 ;
    LAYER V3 ;
    RECT 238.6 140.56 240.6 141.36 ;
    LAYER V3 ;
    RECT 235.48 142.26 237.48 143.06 ;
    LAYER V3 ;
    RECT 238.6 143.96 240.6 144.76 ;
    LAYER V3 ;
    RECT 235.48 145.66 237.48 146.46 ;
    LAYER V3 ;
    RECT 238.6 147.36 240.6 148.16 ;
    LAYER V3 ;
    RECT 235.48 149.06 237.48 149.86 ;
    LAYER V3 ;
    RECT 238.6 150.76 240.6 151.56 ;
    LAYER V3 ;
    RECT 235.48 152.46 237.48 153.26 ;
    LAYER V3 ;
    RECT 238.6 154.16 240.6 154.96 ;
    LAYER V3 ;
    RECT 235.48 155.86 237.48 156.66 ;
    LAYER V3 ;
    RECT 238.6 157.56 240.6 158.36 ;
    LAYER V3 ;
    RECT 235.48 159.26 237.48 160.06 ;
    LAYER V3 ;
    RECT 238.6 160.96 240.6 161.76 ;
    LAYER V3 ;
    RECT 235.48 162.66 237.48 163.46 ;
    LAYER V3 ;
    RECT 238.6 164.36 240.6 165.16 ;
    LAYER V3 ;
    RECT 235.48 166.06 237.48 166.86 ;
    LAYER V3 ;
    RECT 238.6 167.76 240.6 168.56 ;
    LAYER V3 ;
    RECT 235.48 169.46 237.48 170.26 ;
    LAYER V3 ;
    RECT 238.6 171.16 240.6 171.96 ;
    LAYER V3 ;
    RECT 235.48 172.86 237.48 173.66 ;
    LAYER V3 ;
    RECT 238.6 174.56 240.6 175.36 ;
    LAYER V3 ;
    RECT 235.48 176.26 237.48 177.06 ;
    LAYER V3 ;
    RECT 238.6 177.96 240.6 178.76 ;
    LAYER V3 ;
    RECT 235.48 179.66 237.48 180.46 ;
    LAYER V3 ;
    RECT 238.6 181.36 240.6 182.16 ;
    LAYER V3 ;
    RECT 235.48 183.06 237.48 183.86 ;
    LAYER V3 ;
    RECT 238.6 184.76 240.6 185.56 ;
    LAYER V3 ;
    RECT 235.48 186.46 237.48 187.26 ;
    LAYER V3 ;
    RECT 238.6 188.16 240.6 188.96 ;
    LAYER V3 ;
    RECT 235.48 189.86 237.48 190.66 ;
    LAYER V3 ;
    RECT 238.6 191.56 240.6 192.36 ;
    LAYER V3 ;
    RECT 235.48 193.26 237.48 194.06 ;
    LAYER V3 ;
    RECT 238.6 194.96 240.6 195.76 ;
    LAYER V3 ;
    RECT 235.48 196.66 237.48 197.46 ;
    LAYER V3 ;
    RECT 238.6 198.36 240.6 199.16 ;
    LAYER V3 ;
    RECT 235.48 200.06 237.48 200.86 ;
    LAYER V3 ;
    RECT 238.6 201.76 240.6 202.56 ;
    LAYER V3 ;
    RECT 235.48 203.46 237.48 204.26 ;
    LAYER V3 ;
    RECT 238.6 205.16 240.6 205.96 ;
    LAYER V3 ;
    RECT 235.48 206.86 237.48 207.66 ;
    LAYER V3 ;
    RECT 238.6 208.56 240.6 209.36 ;
    LAYER V3 ;
    RECT 235.48 210.26 237.48 211.06 ;
    LAYER V3 ;
    RECT 238.6 211.96 240.6 212.76 ;
    LAYER V3 ;
    RECT 235.48 213.66 237.48 214.46 ;
    LAYER V3 ;
    RECT 238.6 215.36 240.6 216.16 ;
    LAYER V3 ;
    RECT 235.48 217.06 237.48 217.86 ;
    LAYER V3 ;
    RECT 238.6 218.76 240.6 219.56 ;
    LAYER V3 ;
    RECT 235.48 220.46 237.48 221.26 ;
    LAYER V3 ;
    RECT 238.6 222.16 240.6 222.96 ;
    LAYER V3 ;
    RECT 235.48 223.86 237.48 224.66 ;
    LAYER V3 ;
    RECT 238.6 225.56 240.6 226.36 ;
    LAYER V3 ;
    RECT 235.48 227.26 237.48 228.06 ;
    LAYER V3 ;
    RECT 238.6 228.96 240.6 229.76 ;
    LAYER V3 ;
    RECT 235.48 230.66 237.48 231.46 ;
    LAYER V3 ;
    RECT 238.6 232.36 240.6 233.16 ;
    LAYER V3 ;
    RECT 235.48 234.06 237.48 234.86 ;
    LAYER V3 ;
    RECT 238.6 235.76 240.6 236.56 ;
    LAYER V3 ;
    RECT 235.48 237.46 237.48 238.26 ;
    LAYER V3 ;
    RECT 238.6 239.16 240.6 239.96 ;
    LAYER V3 ;
    RECT 235.48 240.86 237.48 241.66 ;
    LAYER V3 ;
    RECT 238.6 242.56 240.6 243.36 ;
    LAYER V3 ;
    RECT 235.48 244.26 237.48 245.06 ;
    LAYER V3 ;
    RECT 238.6 245.96 240.6 246.76 ;
    LAYER V3 ;
    RECT 235.48 247.66 237.48 248.46 ;
    LAYER V3 ;
    RECT 238.6 249.36 240.6 250.16 ;
    LAYER V3 ;
    RECT 235.48 251.06 237.48 251.86 ;
    LAYER V3 ;
    RECT 238.6 252.76 240.6 253.56 ;
    LAYER V3 ;
    RECT 235.48 254.46 237.48 255.26 ;
    LAYER V3 ;
    RECT 238.6 256.16 240.6 256.96 ;
    LAYER V3 ;
    RECT 235.48 257.86 237.48 258.66 ;
    LAYER V3 ;
    RECT 238.6 259.56 240.6 260.36 ;
    LAYER V3 ;
    RECT 235.48 261.26 237.48 262.06 ;
    LAYER V3 ;
    RECT 238.6 262.96 240.6 263.76 ;
    LAYER V3 ;
    RECT 235.48 264.66 237.48 265.46 ;
    LAYER V3 ;
    RECT 238.6 266.36 240.6 267.16 ;
    LAYER V3 ;
    RECT 235.48 268.06 237.48 268.86 ;
    LAYER V3 ;
    RECT 238.6 269.76 240.6 270.56 ;
    LAYER V3 ;
    RECT 235.48 271.46 237.48 272.26 ;
    LAYER V3 ;
    RECT 238.6 273.16 240.6 273.96 ;
    LAYER V3 ;
    RECT 235.48 274.86 237.48 275.66 ;
    LAYER V3 ;
    RECT 238.6 276.56 240.6 277.36 ;
    LAYER V3 ;
    RECT 235.48 278.26 237.48 279.06 ;
    LAYER V3 ;
    RECT 238.6 279.96 240.6 280.76 ;
    LAYER V3 ;
    RECT 235.48 281.66 237.48 282.46 ;
    LAYER V3 ;
    RECT 238.6 283.36 240.6 284.16 ;
    LAYER V3 ;
    RECT 235.48 285.06 237.48 285.86 ;
    LAYER V3 ;
    RECT 238.6 286.76 240.6 287.56 ;
    LAYER V3 ;
    RECT 235.48 288.46 237.48 289.26 ;
    LAYER V3 ;
    RECT 238.6 290.16 240.6 290.96 ;
    LAYER V3 ;
    RECT 235.48 291.86 237.48 292.66 ;
    LAYER V3 ;
    RECT 238.6 293.56 240.6 294.36 ;
    LAYER V3 ;
    RECT 235.48 295.26 237.48 296.06 ;
    LAYER V3 ;
    RECT 238.6 296.96 240.6 297.76 ;
    LAYER V3 ;
    RECT 235.48 298.66 237.48 299.46 ;
    LAYER V3 ;
    RECT 238.6 300.36 240.6 301.16 ;
    LAYER V3 ;
    RECT 235.48 302.06 237.48 302.86 ;
    LAYER V3 ;
    RECT 238.6 303.76 240.6 304.56 ;
    LAYER V3 ;
    RECT 235.48 305.46 237.48 306.26 ;
    LAYER V3 ;
    RECT 238.6 307.16 240.6 307.96 ;
    LAYER V3 ;
    RECT 235.48 308.86 237.48 309.66 ;
    LAYER V3 ;
    RECT 238.6 310.56 240.6 311.36 ;
    LAYER V3 ;
    RECT 235.48 312.26 237.48 313.06 ;
    LAYER V3 ;
    RECT 238.6 313.96 240.6 314.76 ;
    LAYER V3 ;
    RECT 235.48 315.66 237.48 316.46 ;
    LAYER V3 ;
    RECT 238.6 317.36 240.6 318.16 ;
    LAYER V3 ;
    RECT 235.48 319.06 237.48 319.86 ;
    LAYER V3 ;
    RECT 238.6 320.76 240.6 321.56 ;
    LAYER V3 ;
    RECT 235.48 322.46 237.48 323.26 ;
    LAYER V3 ;
    RECT 238.6 324.16 240.6 324.96 ;
    LAYER V3 ;
    RECT 235.48 325.86 237.48 326.66 ;
    LAYER V3 ;
    RECT 238.6 327.56 240.6 328.36 ;
    LAYER V3 ;
    RECT 235.48 329.26 237.48 330.06 ;
    LAYER V3 ;
    RECT 238.6 330.96 240.6 331.76 ;
    LAYER V3 ;
    RECT 235.48 332.66 237.48 333.46 ;
    LAYER V3 ;
    RECT 238.6 334.36 240.6 335.16 ;
    LAYER V3 ;
    RECT 235.48 336.06 237.48 336.86 ;
    LAYER V3 ;
    RECT 238.6 337.76 240.6 338.56 ;
    LAYER V3 ;
    RECT 235.48 339.46 237.48 340.26 ;
    LAYER V3 ;
    RECT 238.6 341.16 240.6 341.96 ;
    LAYER V3 ;
    RECT 235.48 342.86 237.48 343.66 ;
    LAYER V3 ;
    RECT 238.6 344.56 240.6 345.36 ;
    LAYER V3 ;
    RECT 235.48 346.26 237.48 347.06 ;
    LAYER V3 ;
    RECT 238.6 347.96 240.6 348.76 ;
    LAYER V3 ;
    RECT 235.48 349.66 237.48 350.46 ;
    LAYER V3 ;
    RECT 238.6 351.36 240.6 352.16 ;
    LAYER V3 ;
    RECT 235.48 353.06 237.48 353.86 ;
    LAYER V3 ;
    RECT 238.6 354.76 240.6 355.56 ;
    LAYER V3 ;
    RECT 235.48 356.46 237.48 357.26 ;
    LAYER V3 ;
    RECT 238.6 358.16 240.6 358.96 ;
    LAYER V3 ;
    RECT 235.48 359.86 237.48 360.66 ;
    LAYER V3 ;
    RECT 238.6 361.56 240.6 362.36 ;
    LAYER V3 ;
    RECT 235.48 363.26 237.48 364.06 ;
    LAYER V3 ;
    RECT 238.6 364.96 240.6 365.76 ;
    LAYER V3 ;
    RECT 235.48 366.66 237.48 367.46 ;
    LAYER V3 ;
    RECT 238.6 368.36 240.6 369.16 ;
    LAYER V3 ;
    RECT 235.48 370.06 237.48 370.86 ;
    LAYER V3 ;
    RECT 238.6 371.76 240.6 372.56 ;
    LAYER V3 ;
    RECT 235.48 373.46 237.48 374.26 ;
    LAYER V3 ;
    RECT 238.6 375.16 240.6 375.96 ;
    LAYER V3 ;
    RECT 235.48 376.86 237.48 377.66 ;
    LAYER V3 ;
    RECT 238.6 378.56 240.6 379.36 ;
    LAYER V3 ;
    RECT 235.48 380.26 237.48 381.06 ;
    LAYER V3 ;
    RECT 238.6 381.96 240.6 382.76 ;
    LAYER V3 ;
    RECT 235.48 383.66 237.48 384.46 ;
    LAYER V3 ;
    RECT 238.6 385.36 240.6 386.16 ;
    LAYER V3 ;
    RECT 235.48 387.06 237.48 387.86 ;
    LAYER V3 ;
    RECT 238.6 388.76 240.6 389.56 ;
    LAYER V3 ;
    RECT 235.48 390.46 237.48 391.26 ;
    LAYER V3 ;
    RECT 238.6 392.16 240.6 392.96 ;
    LAYER V3 ;
    RECT 235.48 393.86 237.48 394.66 ;
    LAYER V3 ;
    RECT 238.6 395.56 240.6 396.36 ;
    LAYER V3 ;
    RECT 235.48 397.26 237.48 398.06 ;
    LAYER V3 ;
    RECT 238.6 398.96 240.6 399.76 ;
    LAYER V3 ;
    RECT 235.48 400.66 237.48 401.46 ;
    LAYER V3 ;
    RECT 238.6 402.36 240.6 403.16 ;
    LAYER V3 ;
    RECT 235.48 404.06 237.48 404.86 ;
    LAYER V3 ;
    RECT 238.6 405.76 240.6 406.56 ;
    LAYER V3 ;
    RECT 235.48 407.46 237.48 408.26 ;
    LAYER V3 ;
    RECT 238.6 409.16 240.6 409.96 ;
    LAYER V3 ;
    RECT 235.48 410.86 237.48 411.66 ;
    LAYER V3 ;
    RECT 238.6 412.56 240.6 413.36 ;
    LAYER V3 ;
    RECT 235.48 414.26 237.48 415.06 ;
    LAYER V3 ;
    RECT 238.6 415.96 240.6 416.76 ;
    LAYER V3 ;
    RECT 235.48 417.66 237.48 418.46 ;
    LAYER V3 ;
    RECT 238.6 419.36 240.6 420.16 ;
    LAYER V3 ;
    RECT 235.48 421.06 237.48 421.86 ;
    LAYER V3 ;
    RECT 238.6 422.76 240.6 423.56 ;
    LAYER V3 ;
    RECT 235.48 424.46 237.48 425.26 ;
    LAYER V3 ;
    RECT 238.6 426.16 240.6 426.96 ;
    LAYER V3 ;
    RECT 235.48 427.86 237.48 428.66 ;
    LAYER V3 ;
    RECT 238.6 429.56 240.6 430.36 ;
    LAYER V3 ;
    RECT 235.48 431.26 237.48 432.06 ;
    LAYER V3 ;
    RECT 238.6 432.96 240.6 433.76 ;
    LAYER V3 ;
    RECT 235.48 434.66 237.48 435.46 ;
    LAYER V3 ;
    RECT 238.6 436.36 240.6 437.16 ;
    LAYER V3 ;
    RECT 235.48 438.06 237.48 438.86 ;
    LAYER V3 ;
    RECT 238.6 439.76 240.6 440.56 ;
    LAYER V3 ;
    RECT 235.48 441.46 237.48 442.26 ;
    LAYER V3 ;
    RECT 238.6 443.16 240.6 443.96 ;
    LAYER V3 ;
    RECT 235.48 444.86 237.48 445.66 ;
    LAYER V3 ;
    RECT 238.6 446.56 240.6 447.36 ;
    LAYER V3 ;
    RECT 235.48 448.26 237.48 449.06 ;
    LAYER V3 ;
    RECT 238.6 449.96 240.6 450.76 ;
    LAYER V3 ;
    RECT 235.48 451.66 237.48 452.46 ;
    LAYER V3 ;
    RECT 238.6 453.36 240.6 454.16 ;
    LAYER V3 ;
    RECT 235.48 455.06 237.48 455.86 ;
    LAYER V3 ;
    RECT 238.6 456.76 240.6 457.56 ;
    LAYER V3 ;
    RECT 235.48 458.46 237.48 459.26 ;
    LAYER V3 ;
    RECT 238.6 460.16 240.6 460.96 ;
    LAYER V3 ;
    RECT 235.48 461.86 237.48 462.66 ;
    LAYER V3 ;
    RECT 238.6 463.56 240.6 464.36 ;
    LAYER V3 ;
    RECT 235.48 465.26 237.48 466.06 ;
    LAYER V3 ;
    RECT 238.6 466.96 240.6 467.76 ;
    LAYER V3 ;
    RECT 235.48 468.66 237.48 469.46 ;
    LAYER V3 ;
    RECT 238.6 470.36 240.6 471.16 ;
    LAYER V3 ;
    RECT 235.48 472.06 237.48 472.86 ;
    LAYER V3 ;
    RECT 238.6 473.76 240.6 474.56 ;
    LAYER V3 ;
    RECT 235.48 475.46 237.48 476.26 ;
    LAYER V3 ;
    RECT 238.6 477.16 240.6 477.96 ;
    LAYER V3 ;
    RECT 235.48 478.86 237.48 479.66 ;
    LAYER V3 ;
    RECT 238.6 480.56 240.6 481.36 ;
    LAYER V3 ;
    RECT 235.48 482.26 237.48 483.06 ;
    LAYER V3 ;
    RECT 238.6 483.96 240.6 484.76 ;
    LAYER V3 ;
    RECT 235.48 485.66 237.48 486.46 ;
    LAYER V3 ;
    RECT 238.6 487.36 240.6 488.16 ;
    LAYER V3 ;
    RECT 235.48 489.06 237.48 489.86 ;
    LAYER V3 ;
    RECT 238.6 490.76 240.6 491.56 ;
    LAYER V3 ;
    RECT 235.48 492.46 237.48 493.26 ;
    LAYER V3 ;
    RECT 238.6 494.16 240.6 494.96 ;
    LAYER V3 ;
    RECT 235.48 495.86 237.48 496.66 ;
    LAYER V3 ;
    RECT 238.6 497.56 240.6 498.36 ;
    LAYER V3 ;
    RECT 235.48 499.26 237.48 500.06 ;
    LAYER V3 ;
    RECT 238.6 500.96 240.6 501.76 ;
    LAYER V3 ;
    RECT 235.48 502.66 237.48 503.46 ;
    LAYER V3 ;
    RECT 238.6 504.36 240.6 505.16 ;
    LAYER V3 ;
    RECT 238.6 505.6 240.6 506.0 ;
    LAYER V3 ;
    RECT 235.48 506.6 237.48 508.6 ;
    LAYER V3 ;
    RECT 238.6 509.0 240.6 509.8 ;
    LAYER V3 ;
    RECT 0.0 7.94 2.0 9.14 ;
    LAYER V3 ;
    RECT 3.12 12.64 5.12 13.74 ;
    LAYER V3 ;
    RECT 0.0 17.26 2.0 18.46 ;
    LAYER V3 ;
    RECT 3.12 21.41 5.12 22.21 ;
    LAYER V3 ;
    RECT 0.0 25.81 2.0 27.81 ;
    LAYER V3 ;
    RECT 3.12 31.13 5.12 32.13 ;
    LAYER V3 ;
    RECT 3.12 32.98 5.12 33.98 ;
    LAYER V3 ;
    RECT 0.0 35.91 2.0 36.91 ;
    LAYER V3 ;
    RECT 3.12 39.44 5.12 40.44 ;
    LAYER V3 ;
    RECT 3.12 41.29 5.12 42.29 ;
    LAYER V3 ;
    RECT 0.0 50.24 2.0 51.24 ;
    LAYER V3 ;
    RECT 3.12 54.22 5.12 55.22 ;
    LAYER V3 ;
    RECT 0.0 57.02 2.0 58.02 ;
    LAYER V3 ;
    RECT 0.0 60.6 2.0 61.6 ;
    LAYER V3 ;
    RECT 0.0 62.45 2.0 63.45 ;
    LAYER V3 ;
    RECT 0.0 69.16 2.0 69.96 ;
    LAYER V3 ;
    RECT 3.12 70.86 5.12 71.66 ;
    LAYER V3 ;
    RECT 0.0 72.56 2.0 73.36 ;
    LAYER V3 ;
    RECT 3.12 74.26 5.12 75.06 ;
    LAYER V3 ;
    RECT 0.0 75.96 2.0 76.76 ;
    LAYER V3 ;
    RECT 3.12 77.66 5.12 78.46 ;
    LAYER V3 ;
    RECT 0.0 79.36 2.0 80.16 ;
    LAYER V3 ;
    RECT 3.12 81.06 5.12 81.86 ;
    LAYER V3 ;
    RECT 0.0 82.76 2.0 83.56 ;
    LAYER V3 ;
    RECT 3.12 84.46 5.12 85.26 ;
    LAYER V3 ;
    RECT 0.0 86.16 2.0 86.96 ;
    LAYER V3 ;
    RECT 3.12 87.86 5.12 88.66 ;
    LAYER V3 ;
    RECT 0.0 89.56 2.0 90.36 ;
    LAYER V3 ;
    RECT 3.12 91.26 5.12 92.06 ;
    LAYER V3 ;
    RECT 0.0 92.96 2.0 93.76 ;
    LAYER V3 ;
    RECT 3.12 94.66 5.12 95.46 ;
    LAYER V3 ;
    RECT 0.0 96.36 2.0 97.16 ;
    LAYER V3 ;
    RECT 3.12 98.06 5.12 98.86 ;
    LAYER V3 ;
    RECT 0.0 99.76 2.0 100.56 ;
    LAYER V3 ;
    RECT 3.12 101.46 5.12 102.26 ;
    LAYER V3 ;
    RECT 0.0 103.16 2.0 103.96 ;
    LAYER V3 ;
    RECT 3.12 104.86 5.12 105.66 ;
    LAYER V3 ;
    RECT 0.0 106.56 2.0 107.36 ;
    LAYER V3 ;
    RECT 3.12 108.26 5.12 109.06 ;
    LAYER V3 ;
    RECT 0.0 109.96 2.0 110.76 ;
    LAYER V3 ;
    RECT 3.12 111.66 5.12 112.46 ;
    LAYER V3 ;
    RECT 0.0 113.36 2.0 114.16 ;
    LAYER V3 ;
    RECT 3.12 115.06 5.12 115.86 ;
    LAYER V3 ;
    RECT 0.0 116.76 2.0 117.56 ;
    LAYER V3 ;
    RECT 3.12 118.46 5.12 119.26 ;
    LAYER V3 ;
    RECT 0.0 120.16 2.0 120.96 ;
    LAYER V3 ;
    RECT 3.12 121.86 5.12 122.66 ;
    LAYER V3 ;
    RECT 0.0 123.56 2.0 124.36 ;
    LAYER V3 ;
    RECT 3.12 125.26 5.12 126.06 ;
    LAYER V3 ;
    RECT 0.0 126.96 2.0 127.76 ;
    LAYER V3 ;
    RECT 3.12 128.66 5.12 129.46 ;
    LAYER V3 ;
    RECT 0.0 130.36 2.0 131.16 ;
    LAYER V3 ;
    RECT 3.12 132.06 5.12 132.86 ;
    LAYER V3 ;
    RECT 0.0 133.76 2.0 134.56 ;
    LAYER V3 ;
    RECT 3.12 135.46 5.12 136.26 ;
    LAYER V3 ;
    RECT 0.0 137.16 2.0 137.96 ;
    LAYER V3 ;
    RECT 3.12 138.86 5.12 139.66 ;
    LAYER V3 ;
    RECT 0.0 140.56 2.0 141.36 ;
    LAYER V3 ;
    RECT 3.12 142.26 5.12 143.06 ;
    LAYER V3 ;
    RECT 0.0 143.96 2.0 144.76 ;
    LAYER V3 ;
    RECT 3.12 145.66 5.12 146.46 ;
    LAYER V3 ;
    RECT 0.0 147.36 2.0 148.16 ;
    LAYER V3 ;
    RECT 3.12 149.06 5.12 149.86 ;
    LAYER V3 ;
    RECT 0.0 150.76 2.0 151.56 ;
    LAYER V3 ;
    RECT 3.12 152.46 5.12 153.26 ;
    LAYER V3 ;
    RECT 0.0 154.16 2.0 154.96 ;
    LAYER V3 ;
    RECT 3.12 155.86 5.12 156.66 ;
    LAYER V3 ;
    RECT 0.0 157.56 2.0 158.36 ;
    LAYER V3 ;
    RECT 3.12 159.26 5.12 160.06 ;
    LAYER V3 ;
    RECT 0.0 160.96 2.0 161.76 ;
    LAYER V3 ;
    RECT 3.12 162.66 5.12 163.46 ;
    LAYER V3 ;
    RECT 0.0 164.36 2.0 165.16 ;
    LAYER V3 ;
    RECT 3.12 166.06 5.12 166.86 ;
    LAYER V3 ;
    RECT 0.0 167.76 2.0 168.56 ;
    LAYER V3 ;
    RECT 3.12 169.46 5.12 170.26 ;
    LAYER V3 ;
    RECT 0.0 171.16 2.0 171.96 ;
    LAYER V3 ;
    RECT 3.12 172.86 5.12 173.66 ;
    LAYER V3 ;
    RECT 0.0 174.56 2.0 175.36 ;
    LAYER V3 ;
    RECT 3.12 176.26 5.12 177.06 ;
    LAYER V3 ;
    RECT 0.0 177.96 2.0 178.76 ;
    LAYER V3 ;
    RECT 3.12 179.66 5.12 180.46 ;
    LAYER V3 ;
    RECT 0.0 181.36 2.0 182.16 ;
    LAYER V3 ;
    RECT 3.12 183.06 5.12 183.86 ;
    LAYER V3 ;
    RECT 0.0 184.76 2.0 185.56 ;
    LAYER V3 ;
    RECT 3.12 186.46 5.12 187.26 ;
    LAYER V3 ;
    RECT 0.0 188.16 2.0 188.96 ;
    LAYER V3 ;
    RECT 3.12 189.86 5.12 190.66 ;
    LAYER V3 ;
    RECT 0.0 191.56 2.0 192.36 ;
    LAYER V3 ;
    RECT 3.12 193.26 5.12 194.06 ;
    LAYER V3 ;
    RECT 0.0 194.96 2.0 195.76 ;
    LAYER V3 ;
    RECT 3.12 196.66 5.12 197.46 ;
    LAYER V3 ;
    RECT 0.0 198.36 2.0 199.16 ;
    LAYER V3 ;
    RECT 3.12 200.06 5.12 200.86 ;
    LAYER V3 ;
    RECT 0.0 201.76 2.0 202.56 ;
    LAYER V3 ;
    RECT 3.12 203.46 5.12 204.26 ;
    LAYER V3 ;
    RECT 0.0 205.16 2.0 205.96 ;
    LAYER V3 ;
    RECT 3.12 206.86 5.12 207.66 ;
    LAYER V3 ;
    RECT 0.0 208.56 2.0 209.36 ;
    LAYER V3 ;
    RECT 3.12 210.26 5.12 211.06 ;
    LAYER V3 ;
    RECT 0.0 211.96 2.0 212.76 ;
    LAYER V3 ;
    RECT 3.12 213.66 5.12 214.46 ;
    LAYER V3 ;
    RECT 0.0 215.36 2.0 216.16 ;
    LAYER V3 ;
    RECT 3.12 217.06 5.12 217.86 ;
    LAYER V3 ;
    RECT 0.0 218.76 2.0 219.56 ;
    LAYER V3 ;
    RECT 3.12 220.46 5.12 221.26 ;
    LAYER V3 ;
    RECT 0.0 222.16 2.0 222.96 ;
    LAYER V3 ;
    RECT 3.12 223.86 5.12 224.66 ;
    LAYER V3 ;
    RECT 0.0 225.56 2.0 226.36 ;
    LAYER V3 ;
    RECT 3.12 227.26 5.12 228.06 ;
    LAYER V3 ;
    RECT 0.0 228.96 2.0 229.76 ;
    LAYER V3 ;
    RECT 3.12 230.66 5.12 231.46 ;
    LAYER V3 ;
    RECT 0.0 232.36 2.0 233.16 ;
    LAYER V3 ;
    RECT 3.12 234.06 5.12 234.86 ;
    LAYER V3 ;
    RECT 0.0 235.76 2.0 236.56 ;
    LAYER V3 ;
    RECT 3.12 237.46 5.12 238.26 ;
    LAYER V3 ;
    RECT 0.0 239.16 2.0 239.96 ;
    LAYER V3 ;
    RECT 3.12 240.86 5.12 241.66 ;
    LAYER V3 ;
    RECT 0.0 242.56 2.0 243.36 ;
    LAYER V3 ;
    RECT 3.12 244.26 5.12 245.06 ;
    LAYER V3 ;
    RECT 0.0 245.96 2.0 246.76 ;
    LAYER V3 ;
    RECT 3.12 247.66 5.12 248.46 ;
    LAYER V3 ;
    RECT 0.0 249.36 2.0 250.16 ;
    LAYER V3 ;
    RECT 3.12 251.06 5.12 251.86 ;
    LAYER V3 ;
    RECT 0.0 252.76 2.0 253.56 ;
    LAYER V3 ;
    RECT 3.12 254.46 5.12 255.26 ;
    LAYER V3 ;
    RECT 0.0 256.16 2.0 256.96 ;
    LAYER V3 ;
    RECT 3.12 257.86 5.12 258.66 ;
    LAYER V3 ;
    RECT 0.0 259.56 2.0 260.36 ;
    LAYER V3 ;
    RECT 3.12 261.26 5.12 262.06 ;
    LAYER V3 ;
    RECT 0.0 262.96 2.0 263.76 ;
    LAYER V3 ;
    RECT 3.12 264.66 5.12 265.46 ;
    LAYER V3 ;
    RECT 0.0 266.36 2.0 267.16 ;
    LAYER V3 ;
    RECT 3.12 268.06 5.12 268.86 ;
    LAYER V3 ;
    RECT 0.0 269.76 2.0 270.56 ;
    LAYER V3 ;
    RECT 3.12 271.46 5.12 272.26 ;
    LAYER V3 ;
    RECT 0.0 273.16 2.0 273.96 ;
    LAYER V3 ;
    RECT 3.12 274.86 5.12 275.66 ;
    LAYER V3 ;
    RECT 0.0 276.56 2.0 277.36 ;
    LAYER V3 ;
    RECT 3.12 278.26 5.12 279.06 ;
    LAYER V3 ;
    RECT 0.0 279.96 2.0 280.76 ;
    LAYER V3 ;
    RECT 3.12 281.66 5.12 282.46 ;
    LAYER V3 ;
    RECT 0.0 283.36 2.0 284.16 ;
    LAYER V3 ;
    RECT 3.12 285.06 5.12 285.86 ;
    LAYER V3 ;
    RECT 0.0 286.76 2.0 287.56 ;
    LAYER V3 ;
    RECT 3.12 288.46 5.12 289.26 ;
    LAYER V3 ;
    RECT 0.0 290.16 2.0 290.96 ;
    LAYER V3 ;
    RECT 3.12 291.86 5.12 292.66 ;
    LAYER V3 ;
    RECT 0.0 293.56 2.0 294.36 ;
    LAYER V3 ;
    RECT 3.12 295.26 5.12 296.06 ;
    LAYER V3 ;
    RECT 0.0 296.96 2.0 297.76 ;
    LAYER V3 ;
    RECT 3.12 298.66 5.12 299.46 ;
    LAYER V3 ;
    RECT 0.0 300.36 2.0 301.16 ;
    LAYER V3 ;
    RECT 3.12 302.06 5.12 302.86 ;
    LAYER V3 ;
    RECT 0.0 303.76 2.0 304.56 ;
    LAYER V3 ;
    RECT 3.12 305.46 5.12 306.26 ;
    LAYER V3 ;
    RECT 0.0 307.16 2.0 307.96 ;
    LAYER V3 ;
    RECT 3.12 308.86 5.12 309.66 ;
    LAYER V3 ;
    RECT 0.0 310.56 2.0 311.36 ;
    LAYER V3 ;
    RECT 3.12 312.26 5.12 313.06 ;
    LAYER V3 ;
    RECT 0.0 313.96 2.0 314.76 ;
    LAYER V3 ;
    RECT 3.12 315.66 5.12 316.46 ;
    LAYER V3 ;
    RECT 0.0 317.36 2.0 318.16 ;
    LAYER V3 ;
    RECT 3.12 319.06 5.12 319.86 ;
    LAYER V3 ;
    RECT 0.0 320.76 2.0 321.56 ;
    LAYER V3 ;
    RECT 3.12 322.46 5.12 323.26 ;
    LAYER V3 ;
    RECT 0.0 324.16 2.0 324.96 ;
    LAYER V3 ;
    RECT 3.12 325.86 5.12 326.66 ;
    LAYER V3 ;
    RECT 0.0 327.56 2.0 328.36 ;
    LAYER V3 ;
    RECT 3.12 329.26 5.12 330.06 ;
    LAYER V3 ;
    RECT 0.0 330.96 2.0 331.76 ;
    LAYER V3 ;
    RECT 3.12 332.66 5.12 333.46 ;
    LAYER V3 ;
    RECT 0.0 334.36 2.0 335.16 ;
    LAYER V3 ;
    RECT 3.12 336.06 5.12 336.86 ;
    LAYER V3 ;
    RECT 0.0 337.76 2.0 338.56 ;
    LAYER V3 ;
    RECT 3.12 339.46 5.12 340.26 ;
    LAYER V3 ;
    RECT 0.0 341.16 2.0 341.96 ;
    LAYER V3 ;
    RECT 3.12 342.86 5.12 343.66 ;
    LAYER V3 ;
    RECT 0.0 344.56 2.0 345.36 ;
    LAYER V3 ;
    RECT 3.12 346.26 5.12 347.06 ;
    LAYER V3 ;
    RECT 0.0 347.96 2.0 348.76 ;
    LAYER V3 ;
    RECT 3.12 349.66 5.12 350.46 ;
    LAYER V3 ;
    RECT 0.0 351.36 2.0 352.16 ;
    LAYER V3 ;
    RECT 3.12 353.06 5.12 353.86 ;
    LAYER V3 ;
    RECT 0.0 354.76 2.0 355.56 ;
    LAYER V3 ;
    RECT 3.12 356.46 5.12 357.26 ;
    LAYER V3 ;
    RECT 0.0 358.16 2.0 358.96 ;
    LAYER V3 ;
    RECT 3.12 359.86 5.12 360.66 ;
    LAYER V3 ;
    RECT 0.0 361.56 2.0 362.36 ;
    LAYER V3 ;
    RECT 3.12 363.26 5.12 364.06 ;
    LAYER V3 ;
    RECT 0.0 364.96 2.0 365.76 ;
    LAYER V3 ;
    RECT 3.12 366.66 5.12 367.46 ;
    LAYER V3 ;
    RECT 0.0 368.36 2.0 369.16 ;
    LAYER V3 ;
    RECT 3.12 370.06 5.12 370.86 ;
    LAYER V3 ;
    RECT 0.0 371.76 2.0 372.56 ;
    LAYER V3 ;
    RECT 3.12 373.46 5.12 374.26 ;
    LAYER V3 ;
    RECT 0.0 375.16 2.0 375.96 ;
    LAYER V3 ;
    RECT 3.12 376.86 5.12 377.66 ;
    LAYER V3 ;
    RECT 0.0 378.56 2.0 379.36 ;
    LAYER V3 ;
    RECT 3.12 380.26 5.12 381.06 ;
    LAYER V3 ;
    RECT 0.0 381.96 2.0 382.76 ;
    LAYER V3 ;
    RECT 3.12 383.66 5.12 384.46 ;
    LAYER V3 ;
    RECT 0.0 385.36 2.0 386.16 ;
    LAYER V3 ;
    RECT 3.12 387.06 5.12 387.86 ;
    LAYER V3 ;
    RECT 0.0 388.76 2.0 389.56 ;
    LAYER V3 ;
    RECT 3.12 390.46 5.12 391.26 ;
    LAYER V3 ;
    RECT 0.0 392.16 2.0 392.96 ;
    LAYER V3 ;
    RECT 3.12 393.86 5.12 394.66 ;
    LAYER V3 ;
    RECT 0.0 395.56 2.0 396.36 ;
    LAYER V3 ;
    RECT 3.12 397.26 5.12 398.06 ;
    LAYER V3 ;
    RECT 0.0 398.96 2.0 399.76 ;
    LAYER V3 ;
    RECT 3.12 400.66 5.12 401.46 ;
    LAYER V3 ;
    RECT 0.0 402.36 2.0 403.16 ;
    LAYER V3 ;
    RECT 3.12 404.06 5.12 404.86 ;
    LAYER V3 ;
    RECT 0.0 405.76 2.0 406.56 ;
    LAYER V3 ;
    RECT 3.12 407.46 5.12 408.26 ;
    LAYER V3 ;
    RECT 0.0 409.16 2.0 409.96 ;
    LAYER V3 ;
    RECT 3.12 410.86 5.12 411.66 ;
    LAYER V3 ;
    RECT 0.0 412.56 2.0 413.36 ;
    LAYER V3 ;
    RECT 3.12 414.26 5.12 415.06 ;
    LAYER V3 ;
    RECT 0.0 415.96 2.0 416.76 ;
    LAYER V3 ;
    RECT 3.12 417.66 5.12 418.46 ;
    LAYER V3 ;
    RECT 0.0 419.36 2.0 420.16 ;
    LAYER V3 ;
    RECT 3.12 421.06 5.12 421.86 ;
    LAYER V3 ;
    RECT 0.0 422.76 2.0 423.56 ;
    LAYER V3 ;
    RECT 3.12 424.46 5.12 425.26 ;
    LAYER V3 ;
    RECT 0.0 426.16 2.0 426.96 ;
    LAYER V3 ;
    RECT 3.12 427.86 5.12 428.66 ;
    LAYER V3 ;
    RECT 0.0 429.56 2.0 430.36 ;
    LAYER V3 ;
    RECT 3.12 431.26 5.12 432.06 ;
    LAYER V3 ;
    RECT 0.0 432.96 2.0 433.76 ;
    LAYER V3 ;
    RECT 3.12 434.66 5.12 435.46 ;
    LAYER V3 ;
    RECT 0.0 436.36 2.0 437.16 ;
    LAYER V3 ;
    RECT 3.12 438.06 5.12 438.86 ;
    LAYER V3 ;
    RECT 0.0 439.76 2.0 440.56 ;
    LAYER V3 ;
    RECT 3.12 441.46 5.12 442.26 ;
    LAYER V3 ;
    RECT 0.0 443.16 2.0 443.96 ;
    LAYER V3 ;
    RECT 3.12 444.86 5.12 445.66 ;
    LAYER V3 ;
    RECT 0.0 446.56 2.0 447.36 ;
    LAYER V3 ;
    RECT 3.12 448.26 5.12 449.06 ;
    LAYER V3 ;
    RECT 0.0 449.96 2.0 450.76 ;
    LAYER V3 ;
    RECT 3.12 451.66 5.12 452.46 ;
    LAYER V3 ;
    RECT 0.0 453.36 2.0 454.16 ;
    LAYER V3 ;
    RECT 3.12 455.06 5.12 455.86 ;
    LAYER V3 ;
    RECT 0.0 456.76 2.0 457.56 ;
    LAYER V3 ;
    RECT 3.12 458.46 5.12 459.26 ;
    LAYER V3 ;
    RECT 0.0 460.16 2.0 460.96 ;
    LAYER V3 ;
    RECT 3.12 461.86 5.12 462.66 ;
    LAYER V3 ;
    RECT 0.0 463.56 2.0 464.36 ;
    LAYER V3 ;
    RECT 3.12 465.26 5.12 466.06 ;
    LAYER V3 ;
    RECT 0.0 466.96 2.0 467.76 ;
    LAYER V3 ;
    RECT 3.12 468.66 5.12 469.46 ;
    LAYER V3 ;
    RECT 0.0 470.36 2.0 471.16 ;
    LAYER V3 ;
    RECT 3.12 472.06 5.12 472.86 ;
    LAYER V3 ;
    RECT 0.0 473.76 2.0 474.56 ;
    LAYER V3 ;
    RECT 3.12 475.46 5.12 476.26 ;
    LAYER V3 ;
    RECT 0.0 477.16 2.0 477.96 ;
    LAYER V3 ;
    RECT 3.12 478.86 5.12 479.66 ;
    LAYER V3 ;
    RECT 0.0 480.56 2.0 481.36 ;
    LAYER V3 ;
    RECT 3.12 482.26 5.12 483.06 ;
    LAYER V3 ;
    RECT 0.0 483.96 2.0 484.76 ;
    LAYER V3 ;
    RECT 3.12 485.66 5.12 486.46 ;
    LAYER V3 ;
    RECT 0.0 487.36 2.0 488.16 ;
    LAYER V3 ;
    RECT 3.12 489.06 5.12 489.86 ;
    LAYER V3 ;
    RECT 0.0 490.76 2.0 491.56 ;
    LAYER V3 ;
    RECT 3.12 492.46 5.12 493.26 ;
    LAYER V3 ;
    RECT 0.0 494.16 2.0 494.96 ;
    LAYER V3 ;
    RECT 3.12 495.86 5.12 496.66 ;
    LAYER V3 ;
    RECT 0.0 497.56 2.0 498.36 ;
    LAYER V3 ;
    RECT 3.12 499.26 5.12 500.06 ;
    LAYER V3 ;
    RECT 0.0 500.96 2.0 501.76 ;
    LAYER V3 ;
    RECT 3.12 502.66 5.12 503.46 ;
    LAYER V3 ;
    RECT 0.0 504.36 2.0 505.16 ;
    LAYER V3 ;
    RECT 0.0 505.6 2.0 506.0 ;
    LAYER V3 ;
    RECT 3.12 506.6 5.12 508.6 ;
    LAYER V3 ;
    RECT 0.0 509.0 2.0 509.8 ;
    END
  END RA1SHD

END LIBRARY

