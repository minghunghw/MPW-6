VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RA1SHD
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RA1SHD 0 0 ;
  SIZE 240.6 BY 517.18 ;
  SYMMETRY X Y R90 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.45 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.236 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.326 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.525 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 137.81 6.24 138.41 6.84 ;
      LAYER M2 ;
        RECT 137.81 6.24 138.41 6.84 ;
      LAYER M3 ;
        RECT 137.81 6.24 138.41 6.84 ;
      LAYER M4 ;
        RECT 137.81 6.24 138.41 6.84 ;
      LAYER V3 ;
        RECT 138.01 6.44 138.21 6.64 ;
      LAYER V2 ;
        RECT 138.01 6.44 138.21 6.64 ;
      LAYER V1 ;
        RECT 138.01 6.44 138.21 6.64 ;
    END
  END A[0]
  PIN A[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.45 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.236 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.326 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.525 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 93.61 6.24 94.21 6.84 ;
      LAYER M2 ;
        RECT 93.61 6.24 94.21 6.84 ;
      LAYER M3 ;
        RECT 93.61 6.24 94.21 6.84 ;
      LAYER M4 ;
        RECT 93.61 6.24 94.21 6.84 ;
      LAYER V3 ;
        RECT 93.81 6.44 94.01 6.64 ;
      LAYER V2 ;
        RECT 93.81 6.44 94.01 6.64 ;
      LAYER V1 ;
        RECT 93.81 6.44 94.01 6.64 ;
    END
  END A[10]
  PIN A[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.45 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.236 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.326 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.525 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 90.21 6.24 90.81 6.84 ;
      LAYER M2 ;
        RECT 90.21 6.24 90.81 6.84 ;
      LAYER M3 ;
        RECT 90.21 6.24 90.81 6.84 ;
      LAYER M4 ;
        RECT 90.21 6.24 90.81 6.84 ;
      LAYER V3 ;
        RECT 90.41 6.44 90.61 6.64 ;
      LAYER V2 ;
        RECT 90.41 6.44 90.61 6.64 ;
      LAYER V1 ;
        RECT 90.41 6.44 90.61 6.64 ;
    END
  END A[11]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.45 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.236 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.326 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.525 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 134.41 6.24 135.01 6.84 ;
      LAYER M2 ;
        RECT 134.41 6.24 135.01 6.84 ;
      LAYER M3 ;
        RECT 134.41 6.24 135.01 6.84 ;
      LAYER M4 ;
        RECT 134.41 6.24 135.01 6.84 ;
      LAYER V3 ;
        RECT 134.61 6.44 134.81 6.64 ;
      LAYER V2 ;
        RECT 134.61 6.44 134.81 6.64 ;
      LAYER V1 ;
        RECT 134.61 6.44 134.81 6.64 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.45 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.236 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.326 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.525 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 131.01 6.24 131.61 6.84 ;
      LAYER M2 ;
        RECT 131.01 6.24 131.61 6.84 ;
      LAYER M3 ;
        RECT 131.01 6.24 131.61 6.84 ;
      LAYER M4 ;
        RECT 131.01 6.24 131.61 6.84 ;
      LAYER V3 ;
        RECT 131.21 6.44 131.41 6.64 ;
      LAYER V2 ;
        RECT 131.21 6.44 131.41 6.64 ;
      LAYER V1 ;
        RECT 131.21 6.44 131.41 6.64 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.45 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.236 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.326 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.525 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 127.61 6.24 128.21 6.84 ;
      LAYER M2 ;
        RECT 127.61 6.24 128.21 6.84 ;
      LAYER M3 ;
        RECT 127.61 6.24 128.21 6.84 ;
      LAYER M4 ;
        RECT 127.61 6.24 128.21 6.84 ;
      LAYER V3 ;
        RECT 127.81 6.44 128.01 6.64 ;
      LAYER V2 ;
        RECT 127.81 6.44 128.01 6.64 ;
      LAYER V1 ;
        RECT 127.81 6.44 128.01 6.64 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.45 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.236 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.326 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.525 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 120.81 6.24 121.41 6.84 ;
      LAYER M2 ;
        RECT 120.81 6.24 121.41 6.84 ;
      LAYER M3 ;
        RECT 120.81 6.24 121.41 6.84 ;
      LAYER M4 ;
        RECT 120.81 6.24 121.41 6.84 ;
      LAYER V3 ;
        RECT 121.01 6.44 121.21 6.64 ;
      LAYER V2 ;
        RECT 121.01 6.44 121.21 6.64 ;
      LAYER V1 ;
        RECT 121.01 6.44 121.21 6.64 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.45 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.236 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.326 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.525 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 117.41 6.24 118.01 6.84 ;
      LAYER M2 ;
        RECT 117.41 6.24 118.01 6.84 ;
      LAYER M3 ;
        RECT 117.41 6.24 118.01 6.84 ;
      LAYER M4 ;
        RECT 117.41 6.24 118.01 6.84 ;
      LAYER V3 ;
        RECT 117.61 6.44 117.81 6.64 ;
      LAYER V2 ;
        RECT 117.61 6.44 117.81 6.64 ;
      LAYER V1 ;
        RECT 117.61 6.44 117.81 6.64 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.45 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.236 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.326 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.525 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 114.01 6.24 114.61 6.84 ;
      LAYER M2 ;
        RECT 114.01 6.24 114.61 6.84 ;
      LAYER M3 ;
        RECT 114.01 6.24 114.61 6.84 ;
      LAYER M4 ;
        RECT 114.01 6.24 114.61 6.84 ;
      LAYER V3 ;
        RECT 114.21 6.44 114.41 6.64 ;
      LAYER V2 ;
        RECT 114.21 6.44 114.41 6.64 ;
      LAYER V1 ;
        RECT 114.21 6.44 114.41 6.64 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.45 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.236 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.326 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.525 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 107.21 6.24 107.81 6.84 ;
      LAYER M2 ;
        RECT 107.21 6.24 107.81 6.84 ;
      LAYER M3 ;
        RECT 107.21 6.24 107.81 6.84 ;
      LAYER M4 ;
        RECT 107.21 6.24 107.81 6.84 ;
      LAYER V3 ;
        RECT 107.41 6.44 107.61 6.64 ;
      LAYER V2 ;
        RECT 107.41 6.44 107.61 6.64 ;
      LAYER V1 ;
        RECT 107.41 6.44 107.61 6.64 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.45 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.236 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.326 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.525 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 103.81 6.24 104.41 6.84 ;
      LAYER M2 ;
        RECT 103.81 6.24 104.41 6.84 ;
      LAYER M3 ;
        RECT 103.81 6.24 104.41 6.84 ;
      LAYER M4 ;
        RECT 103.81 6.24 104.41 6.84 ;
      LAYER V3 ;
        RECT 104.01 6.44 104.21 6.64 ;
      LAYER V2 ;
        RECT 104.01 6.44 104.21 6.64 ;
      LAYER V1 ;
        RECT 104.01 6.44 104.21 6.64 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.45 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.236 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.326 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.056 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.525 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2112 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 100.41 6.24 101.01 6.84 ;
      LAYER M2 ;
        RECT 100.41 6.24 101.01 6.84 ;
      LAYER M3 ;
        RECT 100.41 6.24 101.01 6.84 ;
      LAYER M4 ;
        RECT 100.41 6.24 101.01 6.84 ;
      LAYER V3 ;
        RECT 100.61 6.44 100.81 6.64 ;
      LAYER V2 ;
        RECT 100.61 6.44 100.81 6.64 ;
      LAYER V1 ;
        RECT 100.61 6.44 100.81 6.64 ;
    END
  END A[9]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.45 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.9 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.65 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.042 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.525 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 144.01 6.24 144.61 6.84 ;
      LAYER M2 ;
        RECT 144.01 6.24 144.61 6.84 ;
      LAYER M3 ;
        RECT 144.01 6.24 144.61 6.84 ;
      LAYER M4 ;
        RECT 144.01 6.24 144.61 6.84 ;
      LAYER V3 ;
        RECT 144.21 6.44 144.41 6.64 ;
      LAYER V2 ;
        RECT 144.21 6.44 144.41 6.64 ;
      LAYER V1 ;
        RECT 144.21 6.44 144.41 6.64 ;
    END
  END CEN
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.322 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 3.78 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.45 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 25.627 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.03 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.525 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.032 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 152.89 6.24 153.49 6.84 ;
      LAYER M2 ;
        RECT 152.89 6.24 153.49 6.84 ;
      LAYER M3 ;
        RECT 152.89 6.24 153.49 6.84 ;
      LAYER M4 ;
        RECT 152.89 6.24 153.49 6.84 ;
      LAYER V3 ;
        RECT 153.09 6.44 153.29 6.64 ;
      LAYER V2 ;
        RECT 153.09 6.44 153.29 6.64 ;
      LAYER V1 ;
        RECT 153.09 6.44 153.29 6.64 ;
    END
  END CLK
  PIN D[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5712 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2848 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 23.71 6.24 24.31 6.84 ;
      LAYER M2 ;
        RECT 23.71 6.24 24.31 6.84 ;
      LAYER M3 ;
        RECT 23.71 6.24 24.31 6.84 ;
      LAYER M4 ;
        RECT 23.71 6.24 24.31 7.04 ;
      LAYER V3 ;
        RECT 23.91 6.44 24.11 6.64 ;
      LAYER V2 ;
        RECT 23.91 6.44 24.11 6.64 ;
      LAYER V1 ;
        RECT 23.91 6.44 24.11 6.64 ;
    END
  END D[0]
  PIN D[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5712 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2848 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 30.91 6.24 31.51 6.84 ;
      LAYER M2 ;
        RECT 30.91 6.24 31.51 6.84 ;
      LAYER M3 ;
        RECT 30.91 6.24 31.51 7.04 ;
      LAYER M4 ;
        RECT 30.91 6.24 31.51 7.04 ;
      LAYER V3 ;
        RECT 31.1 6.44 31.3 6.64 ;
      LAYER V2 ;
        RECT 31.11 6.44 31.31 6.64 ;
      LAYER V1 ;
        RECT 31.11 6.44 31.31 6.64 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5712 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2848 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 63.31 6.24 63.91 6.84 ;
      LAYER M2 ;
        RECT 63.31 6.24 63.91 6.84 ;
      LAYER M3 ;
        RECT 63.31 6.24 63.91 7.04 ;
      LAYER M4 ;
        RECT 63.31 6.24 63.91 7.04 ;
      LAYER V3 ;
        RECT 63.52 6.44 63.72 6.64 ;
      LAYER V2 ;
        RECT 63.51 6.44 63.71 6.64 ;
      LAYER V1 ;
        RECT 63.51 6.44 63.71 6.64 ;
    END
  END D[2]
  PIN D[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5712 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2848 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 70.51 6.24 71.11 6.84 ;
      LAYER M2 ;
        RECT 70.51 6.24 71.11 6.84 ;
      LAYER M3 ;
        RECT 70.51 6.24 71.11 7.04 ;
      LAYER M4 ;
        RECT 70.51 6.24 71.11 7.04 ;
      LAYER V3 ;
        RECT 70.7 6.44 70.9 6.64 ;
      LAYER V2 ;
        RECT 70.71 6.44 70.91 6.64 ;
      LAYER V1 ;
        RECT 70.71 6.44 70.91 6.64 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5712 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2848 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 169.49 6.24 170.09 6.84 ;
      LAYER M2 ;
        RECT 169.49 6.24 170.09 6.84 ;
      LAYER M3 ;
        RECT 169.49 6.24 170.09 7.04 ;
      LAYER M4 ;
        RECT 169.49 6.24 170.09 7.04 ;
      LAYER V3 ;
        RECT 169.7 6.44 169.9 6.64 ;
      LAYER V2 ;
        RECT 169.69 6.44 169.89 6.64 ;
      LAYER V1 ;
        RECT 169.69 6.44 169.89 6.64 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5712 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2848 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 176.69 6.24 177.29 6.84 ;
      LAYER M2 ;
        RECT 176.69 6.24 177.29 6.84 ;
      LAYER M3 ;
        RECT 176.69 6.24 177.29 7.04 ;
      LAYER M4 ;
        RECT 176.69 6.24 177.29 7.04 ;
      LAYER V3 ;
        RECT 176.88 6.44 177.08 6.64 ;
      LAYER V2 ;
        RECT 176.89 6.44 177.09 6.64 ;
      LAYER V1 ;
        RECT 176.89 6.44 177.09 6.64 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5712 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2848 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 209.09 6.24 209.69 6.84 ;
      LAYER M2 ;
        RECT 209.09 6.24 209.69 6.84 ;
      LAYER M3 ;
        RECT 209.09 6.24 209.69 7.04 ;
      LAYER M4 ;
        RECT 209.09 6.24 209.69 7.04 ;
      LAYER V3 ;
        RECT 209.3 6.44 209.5 6.64 ;
      LAYER V2 ;
        RECT 209.29 6.44 209.49 6.64 ;
      LAYER V1 ;
        RECT 209.29 6.44 209.49 6.64 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5712 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2848 LAYER M1 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 216.29 6.24 216.89 6.84 ;
      LAYER M2 ;
        RECT 216.29 6.24 216.89 6.84 ;
      LAYER M3 ;
        RECT 216.29 6.24 216.89 7.04 ;
      LAYER M4 ;
        RECT 216.29 6.24 216.89 7.04 ;
      LAYER V3 ;
        RECT 216.48 6.44 216.68 6.64 ;
      LAYER V2 ;
        RECT 216.49 6.44 216.69 6.64 ;
      LAYER V1 ;
        RECT 216.49 6.44 216.69 6.64 ;
    END
  END D[7]
  PIN Q[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1706 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 1.848 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6208 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 6.468 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 26.11 6.24 26.71 6.84 ;
      LAYER M2 ;
        RECT 26.11 6.24 26.71 6.84 ;
      LAYER M3 ;
        RECT 26.11 6.24 26.71 6.84 ;
      LAYER M4 ;
        RECT 26.11 6.24 26.71 7.04 ;
      LAYER V3 ;
        RECT 26.31 6.44 26.51 6.64 ;
      LAYER V2 ;
        RECT 26.31 6.44 26.51 6.64 ;
      LAYER V1 ;
        RECT 26.31 6.44 26.51 6.64 ;
    END
  END Q[0]
  PIN Q[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1706 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 1.908 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6208 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 6.328 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 28.51 6.24 29.11 6.84 ;
      LAYER M2 ;
        RECT 28.51 6.24 29.11 6.84 ;
      LAYER M3 ;
        RECT 29.01 6.24 29.11 7.04 ;
        RECT 28.51 6.24 29.11 6.84 ;
      LAYER M4 ;
        RECT 28.51 6.24 29.11 7.04 ;
      LAYER V3 ;
        RECT 28.71 6.44 28.91 6.64 ;
      LAYER V2 ;
        RECT 28.71 6.44 28.91 6.64 ;
      LAYER V1 ;
        RECT 28.71 6.44 28.91 6.64 ;
    END
  END Q[1]
  PIN Q[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1706 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 1.908 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6208 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 6.328 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 65.71 6.24 66.31 6.84 ;
      LAYER M2 ;
        RECT 65.71 6.24 66.31 6.84 ;
      LAYER M3 ;
        RECT 65.71 6.24 66.31 6.84 ;
        RECT 65.71 6.24 65.81 7.04 ;
      LAYER M4 ;
        RECT 65.71 6.24 66.31 7.04 ;
      LAYER V3 ;
        RECT 65.91 6.44 66.11 6.64 ;
      LAYER V2 ;
        RECT 65.91 6.44 66.11 6.64 ;
      LAYER V1 ;
        RECT 65.91 6.44 66.11 6.64 ;
    END
  END Q[2]
  PIN Q[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1706 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 1.908 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6208 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 6.328 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 68.11 6.24 68.71 6.84 ;
      LAYER M2 ;
        RECT 68.11 6.24 68.71 6.84 ;
      LAYER M3 ;
        RECT 68.61 6.24 68.71 7.04 ;
        RECT 68.11 6.24 68.71 6.84 ;
      LAYER M4 ;
        RECT 68.11 6.24 68.71 7.04 ;
      LAYER V3 ;
        RECT 68.31 6.44 68.51 6.64 ;
      LAYER V2 ;
        RECT 68.31 6.44 68.51 6.64 ;
      LAYER V1 ;
        RECT 68.31 6.44 68.51 6.64 ;
    END
  END Q[3]
  PIN Q[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1706 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 1.908 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6208 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 6.328 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 171.89 6.24 172.49 6.84 ;
      LAYER M2 ;
        RECT 171.89 6.24 172.49 6.84 ;
      LAYER M3 ;
        RECT 171.89 6.24 172.49 6.84 ;
        RECT 171.89 6.24 171.99 7.04 ;
      LAYER M4 ;
        RECT 171.89 6.24 172.49 7.04 ;
      LAYER V3 ;
        RECT 172.09 6.44 172.29 6.64 ;
      LAYER V2 ;
        RECT 172.09 6.44 172.29 6.64 ;
      LAYER V1 ;
        RECT 172.09 6.44 172.29 6.64 ;
    END
  END Q[4]
  PIN Q[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1706 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 1.908 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6208 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 6.328 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 174.29 6.24 174.89 6.84 ;
      LAYER M2 ;
        RECT 174.29 6.24 174.89 6.84 ;
      LAYER M3 ;
        RECT 174.79 6.24 174.89 7.04 ;
        RECT 174.29 6.24 174.89 6.84 ;
      LAYER M4 ;
        RECT 174.29 6.24 174.89 7.04 ;
      LAYER V3 ;
        RECT 174.49 6.44 174.69 6.64 ;
      LAYER V2 ;
        RECT 174.49 6.44 174.69 6.64 ;
      LAYER V1 ;
        RECT 174.49 6.44 174.69 6.64 ;
    END
  END Q[5]
  PIN Q[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1706 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 1.908 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6208 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 6.328 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 211.49 6.24 212.09 6.84 ;
      LAYER M2 ;
        RECT 211.49 6.24 212.09 6.84 ;
      LAYER M3 ;
        RECT 211.49 6.24 212.09 6.84 ;
        RECT 211.49 6.24 211.59 7.04 ;
      LAYER M4 ;
        RECT 211.49 6.24 212.09 7.04 ;
      LAYER V3 ;
        RECT 211.69 6.44 211.89 6.64 ;
      LAYER V2 ;
        RECT 211.69 6.44 211.89 6.64 ;
      LAYER V1 ;
        RECT 211.69 6.44 211.89 6.64 ;
    END
  END Q[6]
  PIN Q[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1706 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 1.908 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6208 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 6.328 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 213.89 6.24 214.49 6.84 ;
      LAYER M2 ;
        RECT 213.89 6.24 214.49 6.84 ;
      LAYER M3 ;
        RECT 214.39 6.24 214.49 7.04 ;
        RECT 213.89 6.24 214.49 6.84 ;
      LAYER M4 ;
        RECT 213.89 6.24 214.49 7.04 ;
      LAYER V3 ;
        RECT 214.09 6.44 214.29 6.64 ;
      LAYER V2 ;
        RECT 214.09 6.44 214.29 6.64 ;
      LAYER V1 ;
        RECT 214.09 6.44 214.29 6.64 ;
    END
  END Q[7]
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.006 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.97 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.45 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.021 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.535 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.525 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V3 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V1 ;
    PORT
      LAYER M1 ;
        RECT 149.27 6.24 149.87 6.84 ;
      LAYER M2 ;
        RECT 149.27 6.24 149.87 6.84 ;
      LAYER M3 ;
        RECT 149.27 6.24 149.87 6.84 ;
      LAYER M4 ;
        RECT 149.27 6.24 149.87 6.84 ;
      LAYER V3 ;
        RECT 149.47 6.44 149.67 6.64 ;
      LAYER V2 ;
        RECT 149.47 6.44 149.67 6.64 ;
      LAYER V1 ;
        RECT 149.47 6.44 149.67 6.64 ;
    END
  END WEN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M3 ;
        RECT 0 0 1.98 2 ;
    END
    PORT
      LAYER M3 ;
        RECT 238.62 0 240.6 2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M3 ;
        RECT 3.12 3.12 5.1 5.12 ;
    END
    PORT
      LAYER M3 ;
        RECT 235.5 3.12 237.48 5.12 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 232.39 510.04 233.19 510.94 ;
      RECT 231.19 510.04 231.99 510.94 ;
      RECT 227.59 510.04 228.39 510.94 ;
      RECT 226.39 510.04 227.19 510.94 ;
      RECT 222.79 510.04 223.59 510.94 ;
      RECT 221.59 510.04 222.39 510.94 ;
      RECT 217.99 510.04 218.79 510.94 ;
      RECT 216.79 510.04 217.59 510.94 ;
      RECT 213.19 510.04 213.99 510.94 ;
      RECT 211.99 510.04 212.79 510.94 ;
      RECT 208.39 510.04 209.19 510.94 ;
      RECT 207.19 510.04 207.99 510.94 ;
      RECT 203.59 510.04 204.39 510.94 ;
      RECT 202.39 510.04 203.19 510.94 ;
      RECT 198.79 510.04 199.59 510.94 ;
      RECT 197.59 510.04 198.39 510.94 ;
      RECT 193.99 510.04 194.79 510.94 ;
      RECT 192.79 510.04 193.59 510.94 ;
      RECT 191.59 510.04 192.39 510.94 ;
      RECT 187.99 510.04 188.79 510.94 ;
      RECT 186.79 510.04 187.59 510.94 ;
      RECT 183.19 510.04 183.99 510.94 ;
      RECT 181.99 510.04 182.79 510.94 ;
      RECT 178.39 510.04 179.19 510.94 ;
      RECT 177.19 510.04 177.99 510.94 ;
      RECT 173.59 510.04 174.39 510.94 ;
      RECT 172.39 510.04 173.19 510.94 ;
      RECT 168.79 510.04 169.59 510.94 ;
      RECT 167.59 510.04 168.39 510.94 ;
      RECT 163.99 510.04 164.79 510.94 ;
      RECT 162.79 510.04 163.59 510.94 ;
      RECT 159.19 510.04 159.99 510.94 ;
      RECT 157.99 510.04 158.79 510.94 ;
      RECT 154.39 510.04 155.19 510.94 ;
      RECT 153.19 510.04 153.99 510.94 ;
      RECT 150.79 510.04 151.59 510.94 ;
      RECT 149.93 510.04 150.39 510.94 ;
      RECT 231.19 510.04 233.39 510.74 ;
      RECT 226.39 510.04 228.39 510.74 ;
      RECT 221.59 510.04 223.59 510.74 ;
      RECT 216.79 510.04 218.79 510.74 ;
      RECT 211.99 510.04 213.99 510.74 ;
      RECT 207.19 510.04 209.19 510.74 ;
      RECT 202.39 510.04 204.39 510.74 ;
      RECT 197.59 510.04 199.59 510.74 ;
      RECT 191.59 510.04 194.79 510.74 ;
      RECT 186.79 510.04 188.79 510.74 ;
      RECT 181.99 510.04 183.99 510.74 ;
      RECT 177.19 510.04 179.19 510.74 ;
      RECT 172.39 510.04 174.39 510.74 ;
      RECT 167.59 510.04 169.59 510.74 ;
      RECT 162.79 510.04 164.79 510.74 ;
      RECT 157.99 510.04 159.99 510.74 ;
      RECT 153.19 510.04 155.19 510.74 ;
      RECT 153.19 510.04 233.39 510.22 ;
      RECT 149.93 510.04 233.62 510.2 ;
      RECT 233.46 67.81 233.62 510.2 ;
      RECT 231.51 68.88 231.67 510.94 ;
      RECT 230.31 68.88 230.47 510.22 ;
      RECT 229.11 68.88 229.27 510.22 ;
      RECT 227.91 68.88 228.07 510.94 ;
      RECT 226.71 68.88 226.87 510.94 ;
      RECT 225.51 68.88 225.67 510.22 ;
      RECT 224.31 68.88 224.47 510.22 ;
      RECT 223.11 68.88 223.27 510.94 ;
      RECT 221.91 68.88 222.07 510.94 ;
      RECT 220.71 68.88 220.87 510.22 ;
      RECT 219.51 68.88 219.67 510.22 ;
      RECT 218.31 68.88 218.47 510.94 ;
      RECT 217.11 68.88 217.27 510.94 ;
      RECT 215.91 68.88 216.07 510.22 ;
      RECT 214.71 68.88 214.87 510.22 ;
      RECT 213.51 68.88 213.67 510.94 ;
      RECT 212.31 68.88 212.47 510.94 ;
      RECT 211.11 68.88 211.27 510.22 ;
      RECT 209.91 68.88 210.07 510.22 ;
      RECT 208.71 68.88 208.87 510.94 ;
      RECT 207.51 68.88 207.67 510.94 ;
      RECT 206.31 68.88 206.47 510.22 ;
      RECT 205.11 68.88 205.27 510.22 ;
      RECT 203.91 68.88 204.07 510.94 ;
      RECT 202.71 68.88 202.87 510.94 ;
      RECT 201.51 68.88 201.67 510.22 ;
      RECT 200.31 68.88 200.47 510.22 ;
      RECT 199.11 68.88 199.27 510.94 ;
      RECT 197.91 68.88 198.07 510.94 ;
      RECT 196.71 68.88 196.87 510.22 ;
      RECT 195.51 68.88 195.67 510.22 ;
      RECT 194.31 68.88 194.47 510.94 ;
      RECT 191.91 68.88 192.07 510.94 ;
      RECT 190.71 68.88 190.87 510.22 ;
      RECT 189.51 68.88 189.67 510.22 ;
      RECT 188.31 68.88 188.47 510.94 ;
      RECT 187.11 68.88 187.27 510.94 ;
      RECT 185.91 68.88 186.07 510.22 ;
      RECT 184.71 68.88 184.87 510.22 ;
      RECT 183.51 68.88 183.67 510.94 ;
      RECT 182.31 68.88 182.47 510.94 ;
      RECT 181.11 68.88 181.27 510.22 ;
      RECT 179.91 68.88 180.07 510.22 ;
      RECT 178.71 68.88 178.87 510.94 ;
      RECT 177.51 68.88 177.67 510.94 ;
      RECT 176.31 68.88 176.47 510.22 ;
      RECT 175.11 68.88 175.27 510.22 ;
      RECT 173.91 68.88 174.07 510.94 ;
      RECT 172.71 68.88 172.87 510.94 ;
      RECT 171.51 68.88 171.67 510.22 ;
      RECT 170.31 68.88 170.47 510.22 ;
      RECT 169.11 68.88 169.27 510.94 ;
      RECT 167.91 68.88 168.07 510.94 ;
      RECT 166.71 68.88 166.87 510.22 ;
      RECT 165.51 68.88 165.67 510.22 ;
      RECT 164.31 68.88 164.47 510.94 ;
      RECT 163.11 68.88 163.27 510.94 ;
      RECT 161.91 68.88 162.07 510.22 ;
      RECT 160.71 68.88 160.87 510.22 ;
      RECT 159.51 68.88 159.67 510.94 ;
      RECT 158.31 68.88 158.47 510.94 ;
      RECT 157.11 68.88 157.27 510.22 ;
      RECT 155.91 68.88 156.07 510.22 ;
      RECT 154.71 68.88 154.87 510.94 ;
      RECT 152.31 509.46 152.47 510.2 ;
      RECT 153.16 68.88 233.22 509.88 ;
      RECT 152.92 509.46 233.62 509.69 ;
      RECT 152.31 509.46 233.62 509.62 ;
      RECT 152.99 68.88 233.22 509.2 ;
      RECT 233.46 506.6 234.36 508.6 ;
      RECT 150.76 68.88 233.22 505.8 ;
      RECT 149.93 505.2 233.62 505.36 ;
      RECT 233.46 502.66 234.36 503.46 ;
      RECT 233.46 499.26 234.36 500.06 ;
      RECT 233.46 495.86 234.36 496.66 ;
      RECT 233.46 492.46 234.36 493.26 ;
      RECT 233.46 489.06 234.36 489.86 ;
      RECT 233.46 485.66 234.36 486.46 ;
      RECT 233.46 482.26 234.36 483.06 ;
      RECT 233.46 478.86 234.36 479.66 ;
      RECT 233.46 475.46 234.36 476.26 ;
      RECT 233.46 472.06 234.36 472.86 ;
      RECT 233.46 468.66 234.36 469.46 ;
      RECT 233.46 465.26 234.36 466.06 ;
      RECT 233.46 461.86 234.36 462.66 ;
      RECT 233.46 458.46 234.36 459.26 ;
      RECT 233.46 455.06 234.36 455.86 ;
      RECT 233.46 451.66 234.36 452.46 ;
      RECT 233.46 448.26 234.36 449.06 ;
      RECT 233.46 444.86 234.36 445.66 ;
      RECT 233.46 441.46 234.36 442.26 ;
      RECT 233.46 438.06 234.36 438.86 ;
      RECT 233.46 434.66 234.36 435.46 ;
      RECT 233.46 431.26 234.36 432.06 ;
      RECT 233.46 427.86 234.36 428.66 ;
      RECT 233.46 424.46 234.36 425.26 ;
      RECT 233.46 421.06 234.36 421.86 ;
      RECT 233.46 417.66 234.36 418.46 ;
      RECT 233.46 414.26 234.36 415.06 ;
      RECT 233.46 410.86 234.36 411.66 ;
      RECT 233.46 407.46 234.36 408.26 ;
      RECT 233.46 404.06 234.36 404.86 ;
      RECT 233.46 400.66 234.36 401.46 ;
      RECT 233.46 397.26 234.36 398.06 ;
      RECT 233.46 393.86 234.36 394.66 ;
      RECT 233.46 390.46 234.36 391.26 ;
      RECT 233.46 387.06 234.36 387.86 ;
      RECT 233.46 383.66 234.36 384.46 ;
      RECT 233.46 380.26 234.36 381.06 ;
      RECT 233.46 376.86 234.36 377.66 ;
      RECT 233.46 373.46 234.36 374.26 ;
      RECT 233.46 370.06 234.36 370.86 ;
      RECT 233.46 366.66 234.36 367.46 ;
      RECT 233.46 363.26 234.36 364.06 ;
      RECT 233.46 359.86 234.36 360.66 ;
      RECT 233.46 356.46 234.36 357.26 ;
      RECT 233.46 353.06 234.36 353.86 ;
      RECT 233.46 349.66 234.36 350.46 ;
      RECT 233.46 346.26 234.36 347.06 ;
      RECT 233.46 342.86 234.36 343.66 ;
      RECT 233.46 339.46 234.36 340.26 ;
      RECT 233.46 336.06 234.36 336.86 ;
      RECT 233.46 332.66 234.36 333.46 ;
      RECT 233.46 329.26 234.36 330.06 ;
      RECT 233.46 325.86 234.36 326.66 ;
      RECT 233.46 322.46 234.36 323.26 ;
      RECT 233.46 319.06 234.36 319.86 ;
      RECT 233.46 315.66 234.36 316.46 ;
      RECT 233.46 312.26 234.36 313.06 ;
      RECT 233.46 308.86 234.36 309.66 ;
      RECT 233.46 305.46 234.36 306.26 ;
      RECT 233.46 302.06 234.36 302.86 ;
      RECT 233.46 298.66 234.36 299.46 ;
      RECT 233.46 295.26 234.36 296.06 ;
      RECT 233.46 291.86 234.36 292.66 ;
      RECT 233.46 288.46 234.36 289.26 ;
      RECT 233.46 285.06 234.36 285.86 ;
      RECT 233.46 281.66 234.36 282.46 ;
      RECT 233.46 278.26 234.36 279.06 ;
      RECT 233.46 274.86 234.36 275.66 ;
      RECT 233.46 271.46 234.36 272.26 ;
      RECT 233.46 268.06 234.36 268.86 ;
      RECT 233.46 264.66 234.36 265.46 ;
      RECT 233.46 261.26 234.36 262.06 ;
      RECT 233.46 257.86 234.36 258.66 ;
      RECT 233.46 254.46 234.36 255.26 ;
      RECT 233.46 251.06 234.36 251.86 ;
      RECT 233.46 247.66 234.36 248.46 ;
      RECT 233.46 244.26 234.36 245.06 ;
      RECT 233.46 240.86 234.36 241.66 ;
      RECT 233.46 237.46 234.36 238.26 ;
      RECT 233.46 234.06 234.36 234.86 ;
      RECT 233.46 230.66 234.36 231.46 ;
      RECT 233.46 227.26 234.36 228.06 ;
      RECT 233.46 223.86 234.36 224.66 ;
      RECT 233.46 220.46 234.36 221.26 ;
      RECT 233.46 217.06 234.36 217.86 ;
      RECT 233.46 213.66 234.36 214.46 ;
      RECT 233.46 210.26 234.36 211.06 ;
      RECT 233.46 206.86 234.36 207.66 ;
      RECT 233.46 203.46 234.36 204.26 ;
      RECT 233.46 200.06 234.36 200.86 ;
      RECT 233.46 196.66 234.36 197.46 ;
      RECT 233.46 193.26 234.36 194.06 ;
      RECT 233.46 189.86 234.36 190.66 ;
      RECT 233.46 186.46 234.36 187.26 ;
      RECT 233.46 183.06 234.36 183.86 ;
      RECT 233.46 179.66 234.36 180.46 ;
      RECT 233.46 176.26 234.36 177.06 ;
      RECT 233.46 172.86 234.36 173.66 ;
      RECT 233.46 169.46 234.36 170.26 ;
      RECT 233.46 166.06 234.36 166.86 ;
      RECT 233.46 162.66 234.36 163.46 ;
      RECT 233.46 159.26 234.36 160.06 ;
      RECT 233.46 155.86 234.36 156.66 ;
      RECT 233.46 152.46 234.36 153.26 ;
      RECT 233.46 149.06 234.36 149.86 ;
      RECT 233.46 145.66 234.36 146.46 ;
      RECT 233.46 142.26 234.36 143.06 ;
      RECT 233.46 138.86 234.36 139.66 ;
      RECT 233.46 135.46 234.36 136.26 ;
      RECT 233.46 132.06 234.36 132.86 ;
      RECT 233.46 128.66 234.36 129.46 ;
      RECT 233.46 125.26 234.36 126.06 ;
      RECT 233.46 121.86 234.36 122.66 ;
      RECT 233.46 118.46 234.36 119.26 ;
      RECT 233.46 115.06 234.36 115.86 ;
      RECT 233.46 111.66 234.36 112.46 ;
      RECT 233.46 108.26 234.36 109.06 ;
      RECT 233.46 104.86 234.36 105.66 ;
      RECT 233.46 101.46 234.36 102.26 ;
      RECT 233.46 98.06 234.36 98.86 ;
      RECT 233.46 94.66 234.36 95.46 ;
      RECT 233.46 91.26 234.36 92.06 ;
      RECT 233.46 87.86 234.36 88.66 ;
      RECT 233.46 84.46 234.36 85.26 ;
      RECT 233.46 81.06 234.36 81.86 ;
      RECT 233.46 77.66 234.36 78.46 ;
      RECT 233.46 74.26 234.36 75.06 ;
      RECT 233.46 70.86 234.36 71.66 ;
      RECT 149.71 69.07 233.62 69.3 ;
      RECT 149.71 68.83 150.31 69.3 ;
      RECT 233.14 67.81 233.62 68.09 ;
      RECT 233.14 8.2 233.36 68.09 ;
      RECT 233.14 54.22 234.36 55.22 ;
      RECT 233.14 41.29 234.36 42.29 ;
      RECT 233.14 39.44 234.36 40.44 ;
      RECT 233.14 32.98 234.36 33.98 ;
      RECT 233.14 31.13 234.36 32.13 ;
      RECT 233.14 21.41 234.36 22.21 ;
      RECT 233.14 12.64 234.36 13.74 ;
      RECT 232.11 46.75 232.27 47.43 ;
      RECT 231.79 46.75 232.27 46.91 ;
      RECT 231.79 44.23 231.95 46.91 ;
      RECT 154.11 68.47 232.27 68.63 ;
      RECT 232.11 56.96 232.27 68.63 ;
      RECT 229.71 56.96 229.87 68.63 ;
      RECT 227.31 56.96 227.47 68.63 ;
      RECT 224.91 56.96 225.07 68.63 ;
      RECT 222.51 56.96 222.67 68.63 ;
      RECT 220.11 56.96 220.27 68.63 ;
      RECT 217.71 56.96 217.87 68.63 ;
      RECT 215.31 56.96 215.47 68.63 ;
      RECT 212.91 56.96 213.07 68.63 ;
      RECT 210.51 56.96 210.67 68.63 ;
      RECT 208.11 56.96 208.27 68.63 ;
      RECT 205.71 56.96 205.87 68.63 ;
      RECT 203.31 56.96 203.47 68.63 ;
      RECT 200.91 56.96 201.07 68.63 ;
      RECT 198.51 56.96 198.67 68.63 ;
      RECT 196.11 56.96 196.27 68.63 ;
      RECT 193.71 56.96 193.87 68.63 ;
      RECT 192.51 56.96 192.67 68.63 ;
      RECT 190.11 56.96 190.27 68.63 ;
      RECT 187.71 56.96 187.87 68.63 ;
      RECT 185.31 56.96 185.47 68.63 ;
      RECT 182.91 56.96 183.07 68.63 ;
      RECT 180.51 56.96 180.67 68.63 ;
      RECT 178.11 56.96 178.27 68.63 ;
      RECT 175.71 56.96 175.87 68.63 ;
      RECT 173.31 56.96 173.47 68.63 ;
      RECT 170.91 56.96 171.07 68.63 ;
      RECT 168.51 56.96 168.67 68.63 ;
      RECT 166.11 56.96 166.27 68.63 ;
      RECT 163.71 56.96 163.87 68.63 ;
      RECT 161.31 56.96 161.47 68.63 ;
      RECT 158.91 56.96 159.07 68.63 ;
      RECT 156.51 56.96 156.67 68.63 ;
      RECT 154.11 56.96 154.27 68.63 ;
      RECT 229.89 34.88 232.09 35.04 ;
      RECT 231.81 34.59 232.09 35.04 ;
      RECT 230.87 34.59 231.11 35.04 ;
      RECT 229.89 34.59 230.17 35.04 ;
      RECT 230.87 38.38 231.11 39.02 ;
      RECT 231.81 38.38 232.09 38.83 ;
      RECT 229.89 38.38 230.17 38.83 ;
      RECT 229.89 38.38 232.09 38.54 ;
      RECT 230.05 36.47 231.93 36.63 ;
      RECT 231.77 35.88 231.93 36.63 ;
      RECT 230.91 35.23 231.07 36.63 ;
      RECT 230.05 35.88 230.21 36.63 ;
      RECT 231.87 35.23 232.03 36.06 ;
      RECT 229.95 35.23 230.11 36.06 ;
      RECT 231.87 37.11 232.03 38.19 ;
      RECT 230.91 36.79 231.07 38.19 ;
      RECT 229.95 37.11 230.11 38.19 ;
      RECT 231.77 36.79 231.93 37.39 ;
      RECT 230.05 36.79 230.21 37.39 ;
      RECT 230.05 36.79 231.93 36.95 ;
      RECT 230.13 68.07 231.95 68.23 ;
      RECT 230.13 62.02 230.29 68.23 ;
      RECT 230.13 62.02 230.51 62.18 ;
      RECT 230.35 57.45 230.51 62.18 ;
      RECT 230.35 57.45 231.95 57.61 ;
      RECT 231.63 57.39 231.95 57.61 ;
      RECT 231.63 53.74 231.79 57.61 ;
      RECT 231.79 51.32 231.95 53.9 ;
      RECT 231.47 51.32 231.95 51.48 ;
      RECT 231.47 49.88 231.63 51.48 ;
      RECT 231.15 49.88 231.63 50.04 ;
      RECT 231.15 47.71 231.31 50.04 ;
      RECT 230.69 47.71 231.31 47.99 ;
      RECT 231.47 47.39 231.63 49.72 ;
      RECT 231.15 47.39 231.63 47.55 ;
      RECT 231.15 43.85 231.31 47.55 ;
      RECT 231.15 43.85 231.93 44.01 ;
      RECT 231.77 39.56 231.93 44.01 ;
      RECT 231.59 39.56 231.93 39.84 ;
      RECT 231.59 39.16 231.75 39.84 ;
      RECT 231.63 62.9 231.79 67.89 ;
      RECT 231.51 64.59 231.79 65.31 ;
      RECT 230.87 52.58 231.63 52.86 ;
      RECT 231.47 51.64 231.63 52.86 ;
      RECT 230.87 52.18 231.03 52.86 ;
      RECT 231.27 34.44 231.61 34.72 ;
      RECT 231.27 32.44 231.43 34.72 ;
      RECT 231.27 33.11 231.61 33.39 ;
      RECT 231.27 32.44 231.61 32.72 ;
      RECT 231.27 40.7 231.61 40.98 ;
      RECT 231.27 38.7 231.43 40.98 ;
      RECT 231.27 40.03 231.61 40.31 ;
      RECT 231.27 38.7 231.61 38.98 ;
      RECT 231.33 53.23 231.61 53.51 ;
      RECT 231.33 53.03 231.49 53.51 ;
      RECT 230.51 53.03 231.49 53.19 ;
      RECT 230.51 50.98 230.67 53.19 ;
      RECT 230.47 52.54 230.67 52.82 ;
      RECT 230.13 50.98 230.67 51.14 ;
      RECT 230.13 50.8 230.35 51.14 ;
      RECT 230.03 56.67 230.19 61.86 ;
      RECT 230.03 56.67 231.47 56.83 ;
      RECT 231.31 56 231.47 56.83 ;
      RECT 230.19 54.4 230.35 56.83 ;
      RECT 223.47 12.95 231.31 13.55 ;
      RECT 230.71 8.34 231.31 13.55 ;
      RECT 223.47 8.34 224.07 13.55 ;
      RECT 223.47 8.34 231.31 8.88 ;
      RECT 223.47 26.87 231.31 27.47 ;
      RECT 230.71 18.71 231.31 27.47 ;
      RECT 223.47 18.71 224.07 27.47 ;
      RECT 223.47 24.41 231.31 25.01 ;
      RECT 223.47 18.71 231.31 19.31 ;
      RECT 231.15 50.66 231.31 51.5 ;
      RECT 230.51 50.66 231.31 50.82 ;
      RECT 230.51 50.18 230.67 50.82 ;
      RECT 230.03 50.18 230.67 50.5 ;
      RECT 230.03 47.07 230.19 50.5 ;
      RECT 230.03 47.07 230.51 47.23 ;
      RECT 230.35 45.44 230.51 47.23 ;
      RECT 230.91 55.68 231.07 56.51 ;
      RECT 230.91 55.68 231.31 55.84 ;
      RECT 231.15 53.67 231.31 55.84 ;
      RECT 230.67 53.67 231.31 53.83 ;
      RECT 230.67 53.35 230.95 53.83 ;
      RECT 231.15 62.9 231.31 67.89 ;
      RECT 231.09 65.82 231.31 66.55 ;
      RECT 230.83 51.7 231.21 51.92 ;
      RECT 230.83 50.98 230.99 51.92 ;
      RECT 230.35 47.39 230.51 49.72 ;
      RECT 230.35 47.39 230.83 47.55 ;
      RECT 230.67 43.85 230.83 47.55 ;
      RECT 230.05 43.85 230.83 44.01 ;
      RECT 230.05 39.56 230.21 44.01 ;
      RECT 230.05 39.56 230.39 39.84 ;
      RECT 230.23 39.16 230.39 39.84 ;
      RECT 230.37 34.44 230.71 34.72 ;
      RECT 230.55 32.44 230.71 34.72 ;
      RECT 230.37 33.11 230.71 33.39 ;
      RECT 230.37 32.44 230.71 32.72 ;
      RECT 230.37 40.7 230.71 40.98 ;
      RECT 230.55 38.7 230.71 40.98 ;
      RECT 230.37 40.03 230.71 40.31 ;
      RECT 230.37 38.7 230.71 38.98 ;
      RECT 230.51 54.06 230.67 56.51 ;
      RECT 230.15 54.06 230.67 54.22 ;
      RECT 230.15 52.98 230.35 54.22 ;
      RECT 230.15 51.34 230.31 54.22 ;
      RECT 230.15 51.34 230.35 52.12 ;
      RECT 229.71 46.75 229.87 47.43 ;
      RECT 229.39 46.75 230.19 46.91 ;
      RECT 230.03 44.23 230.19 46.91 ;
      RECT 229.39 44.23 229.55 46.91 ;
      RECT 227.49 34.88 229.69 35.04 ;
      RECT 229.41 34.59 229.69 35.04 ;
      RECT 228.47 34.59 228.71 35.04 ;
      RECT 227.49 34.59 227.77 35.04 ;
      RECT 228.47 38.38 228.71 39.02 ;
      RECT 229.41 38.38 229.69 38.83 ;
      RECT 227.49 38.38 227.77 38.83 ;
      RECT 227.49 38.38 229.69 38.54 ;
      RECT 227.65 36.47 229.53 36.63 ;
      RECT 229.37 35.86 229.53 36.63 ;
      RECT 228.51 35.23 228.67 36.63 ;
      RECT 227.65 35.86 227.81 36.63 ;
      RECT 229.47 35.23 229.63 36.05 ;
      RECT 227.55 35.23 227.71 36.05 ;
      RECT 229.47 37.11 229.63 38.19 ;
      RECT 228.51 36.79 228.67 38.19 ;
      RECT 227.55 37.11 227.71 38.19 ;
      RECT 229.37 36.79 229.53 37.39 ;
      RECT 227.65 36.79 227.81 37.39 ;
      RECT 227.65 36.79 229.53 36.95 ;
      RECT 228.27 50.66 228.43 51.5 ;
      RECT 228.27 50.66 229.07 50.82 ;
      RECT 228.91 50.18 229.07 50.82 ;
      RECT 228.91 50.18 229.55 50.5 ;
      RECT 229.39 47.07 229.55 50.5 ;
      RECT 229.07 47.07 229.55 47.23 ;
      RECT 229.07 45.44 229.23 47.23 ;
      RECT 229.39 56.67 229.55 61.86 ;
      RECT 228.11 56.67 229.55 56.83 ;
      RECT 229.23 54.4 229.39 56.83 ;
      RECT 228.11 56 228.27 56.83 ;
      RECT 229.07 47.39 229.23 49.72 ;
      RECT 228.75 47.39 229.23 47.55 ;
      RECT 228.75 43.85 228.91 47.55 ;
      RECT 228.75 43.85 229.53 44.01 ;
      RECT 229.37 39.56 229.53 44.01 ;
      RECT 229.19 39.56 229.53 39.84 ;
      RECT 229.19 39.16 229.35 39.84 ;
      RECT 227.97 53.23 228.25 53.51 ;
      RECT 228.09 53.03 228.25 53.51 ;
      RECT 228.09 53.03 229.07 53.19 ;
      RECT 228.91 50.98 229.07 53.19 ;
      RECT 228.91 52.54 229.11 52.82 ;
      RECT 228.91 50.98 229.45 51.14 ;
      RECT 229.23 50.8 229.45 51.14 ;
      RECT 227.63 68.07 229.45 68.23 ;
      RECT 229.29 62.02 229.45 68.23 ;
      RECT 229.07 62.02 229.45 62.18 ;
      RECT 229.07 57.45 229.23 62.18 ;
      RECT 227.63 57.45 229.23 57.61 ;
      RECT 227.63 57.39 227.95 57.61 ;
      RECT 227.79 53.74 227.95 57.61 ;
      RECT 227.63 51.32 227.79 53.9 ;
      RECT 227.63 51.32 228.11 51.48 ;
      RECT 227.95 49.88 228.11 51.48 ;
      RECT 227.95 49.88 228.43 50.04 ;
      RECT 228.27 47.71 228.43 50.04 ;
      RECT 228.27 47.71 228.89 47.99 ;
      RECT 228.91 54.06 229.07 56.51 ;
      RECT 228.91 54.06 229.43 54.22 ;
      RECT 229.27 51.34 229.43 54.22 ;
      RECT 229.23 52.98 229.43 54.22 ;
      RECT 229.23 51.34 229.43 52.12 ;
      RECT 228.87 34.44 229.21 34.72 ;
      RECT 228.87 32.44 229.03 34.72 ;
      RECT 228.87 33.11 229.21 33.39 ;
      RECT 228.87 32.44 229.21 32.72 ;
      RECT 228.87 40.7 229.21 40.98 ;
      RECT 228.87 38.7 229.03 40.98 ;
      RECT 228.87 40.03 229.21 40.31 ;
      RECT 228.87 38.7 229.21 38.98 ;
      RECT 228.51 55.68 228.67 56.51 ;
      RECT 228.27 55.68 228.67 55.84 ;
      RECT 228.27 53.67 228.43 55.84 ;
      RECT 228.27 53.67 228.91 53.83 ;
      RECT 228.63 53.35 228.91 53.83 ;
      RECT 228.37 51.7 228.75 51.92 ;
      RECT 228.59 50.98 228.75 51.92 ;
      RECT 227.95 52.58 228.71 52.86 ;
      RECT 228.55 52.18 228.71 52.86 ;
      RECT 227.95 51.64 228.11 52.86 ;
      RECT 228.27 62.9 228.43 67.89 ;
      RECT 228.27 65.82 228.49 66.55 ;
      RECT 227.95 47.39 228.11 49.72 ;
      RECT 227.95 47.39 228.43 47.55 ;
      RECT 228.27 43.85 228.43 47.55 ;
      RECT 227.65 43.85 228.43 44.01 ;
      RECT 227.65 39.56 227.81 44.01 ;
      RECT 227.65 39.56 227.99 39.84 ;
      RECT 227.83 39.16 227.99 39.84 ;
      RECT 227.97 34.44 228.31 34.72 ;
      RECT 228.15 32.44 228.31 34.72 ;
      RECT 227.97 33.11 228.31 33.39 ;
      RECT 227.97 32.44 228.31 32.72 ;
      RECT 227.97 40.7 228.31 40.98 ;
      RECT 228.15 38.7 228.31 40.98 ;
      RECT 227.97 40.03 228.31 40.31 ;
      RECT 227.97 38.7 228.31 38.98 ;
      RECT 227.79 62.9 227.95 67.89 ;
      RECT 227.79 64.59 228.07 65.31 ;
      RECT 227.31 46.75 227.47 47.43 ;
      RECT 226.99 46.75 227.79 46.91 ;
      RECT 227.63 44.23 227.79 46.91 ;
      RECT 226.99 44.23 227.15 46.91 ;
      RECT 225.09 34.88 227.29 35.04 ;
      RECT 227.01 34.59 227.29 35.04 ;
      RECT 226.07 34.59 226.31 35.04 ;
      RECT 225.09 34.59 225.37 35.04 ;
      RECT 226.07 38.38 226.31 39.02 ;
      RECT 227.01 38.38 227.29 38.83 ;
      RECT 225.09 38.38 225.37 38.83 ;
      RECT 225.09 38.38 227.29 38.54 ;
      RECT 225.25 36.47 227.13 36.63 ;
      RECT 226.97 35.88 227.13 36.63 ;
      RECT 226.11 35.23 226.27 36.63 ;
      RECT 225.25 35.88 225.41 36.63 ;
      RECT 227.07 35.23 227.23 36.06 ;
      RECT 225.15 35.23 225.31 36.06 ;
      RECT 227.07 37.11 227.23 38.19 ;
      RECT 226.11 36.79 226.27 38.19 ;
      RECT 225.15 37.11 225.31 38.19 ;
      RECT 226.97 36.79 227.13 37.39 ;
      RECT 225.25 36.79 225.41 37.39 ;
      RECT 225.25 36.79 227.13 36.95 ;
      RECT 225.33 68.07 227.15 68.23 ;
      RECT 225.33 62.02 225.49 68.23 ;
      RECT 225.33 62.02 225.71 62.18 ;
      RECT 225.55 57.45 225.71 62.18 ;
      RECT 225.55 57.45 227.15 57.61 ;
      RECT 226.83 57.39 227.15 57.61 ;
      RECT 226.83 53.74 226.99 57.61 ;
      RECT 226.99 51.32 227.15 53.9 ;
      RECT 226.67 51.32 227.15 51.48 ;
      RECT 226.67 49.88 226.83 51.48 ;
      RECT 226.35 49.88 226.83 50.04 ;
      RECT 226.35 47.71 226.51 50.04 ;
      RECT 225.89 47.71 226.51 47.99 ;
      RECT 226.67 47.39 226.83 49.72 ;
      RECT 226.35 47.39 226.83 47.55 ;
      RECT 226.35 43.85 226.51 47.55 ;
      RECT 226.35 43.85 227.13 44.01 ;
      RECT 226.97 39.56 227.13 44.01 ;
      RECT 226.79 39.56 227.13 39.84 ;
      RECT 226.79 39.16 226.95 39.84 ;
      RECT 226.83 62.9 226.99 67.89 ;
      RECT 226.71 64.59 226.99 65.31 ;
      RECT 226.07 52.58 226.83 52.86 ;
      RECT 226.67 51.64 226.83 52.86 ;
      RECT 226.07 52.18 226.23 52.86 ;
      RECT 226.47 34.44 226.81 34.72 ;
      RECT 226.47 32.44 226.63 34.72 ;
      RECT 226.47 33.11 226.81 33.39 ;
      RECT 226.47 32.44 226.81 32.72 ;
      RECT 226.47 40.7 226.81 40.98 ;
      RECT 226.47 38.7 226.63 40.98 ;
      RECT 226.47 40.03 226.81 40.31 ;
      RECT 226.47 38.7 226.81 38.98 ;
      RECT 226.53 53.23 226.81 53.51 ;
      RECT 226.53 53.03 226.69 53.51 ;
      RECT 225.71 53.03 226.69 53.19 ;
      RECT 225.71 50.98 225.87 53.19 ;
      RECT 225.67 52.54 225.87 52.82 ;
      RECT 225.33 50.98 225.87 51.14 ;
      RECT 225.33 50.8 225.55 51.14 ;
      RECT 225.23 56.67 225.39 61.86 ;
      RECT 225.23 56.67 226.67 56.83 ;
      RECT 226.51 56 226.67 56.83 ;
      RECT 225.39 54.4 225.55 56.83 ;
      RECT 226.35 50.66 226.51 51.5 ;
      RECT 225.71 50.66 226.51 50.82 ;
      RECT 225.71 50.18 225.87 50.82 ;
      RECT 225.23 50.18 225.87 50.5 ;
      RECT 225.23 47.07 225.39 50.5 ;
      RECT 225.23 47.07 225.71 47.23 ;
      RECT 225.55 45.44 225.71 47.23 ;
      RECT 226.11 55.68 226.27 56.51 ;
      RECT 226.11 55.68 226.51 55.84 ;
      RECT 226.35 53.67 226.51 55.84 ;
      RECT 225.87 53.67 226.51 53.83 ;
      RECT 225.87 53.35 226.15 53.83 ;
      RECT 226.35 62.9 226.51 67.89 ;
      RECT 226.29 65.82 226.51 66.55 ;
      RECT 226.03 51.7 226.41 51.92 ;
      RECT 226.03 50.98 226.19 51.92 ;
      RECT 225.55 47.39 225.71 49.72 ;
      RECT 225.55 47.39 226.03 47.55 ;
      RECT 225.87 43.85 226.03 47.55 ;
      RECT 225.25 43.85 226.03 44.01 ;
      RECT 225.25 39.56 225.41 44.01 ;
      RECT 225.25 39.56 225.59 39.84 ;
      RECT 225.43 39.16 225.59 39.84 ;
      RECT 225.57 34.44 225.91 34.72 ;
      RECT 225.75 32.44 225.91 34.72 ;
      RECT 225.57 33.11 225.91 33.39 ;
      RECT 225.57 32.44 225.91 32.72 ;
      RECT 225.57 40.7 225.91 40.98 ;
      RECT 225.75 38.7 225.91 40.98 ;
      RECT 225.57 40.03 225.91 40.31 ;
      RECT 225.57 38.7 225.91 38.98 ;
      RECT 225.71 54.06 225.87 56.51 ;
      RECT 225.35 54.06 225.87 54.22 ;
      RECT 225.35 52.98 225.55 54.22 ;
      RECT 225.35 51.34 225.51 54.22 ;
      RECT 225.35 51.34 225.55 52.12 ;
      RECT 224.91 46.75 225.07 47.43 ;
      RECT 224.59 46.75 225.39 46.91 ;
      RECT 225.23 44.23 225.39 46.91 ;
      RECT 224.59 44.23 224.75 46.91 ;
      RECT 222.69 34.88 224.89 35.04 ;
      RECT 224.61 34.59 224.89 35.04 ;
      RECT 223.67 34.59 223.91 35.04 ;
      RECT 222.69 34.59 222.97 35.04 ;
      RECT 223.67 38.38 223.91 39.02 ;
      RECT 224.61 38.38 224.89 38.83 ;
      RECT 222.69 38.38 222.97 38.83 ;
      RECT 222.69 38.38 224.89 38.54 ;
      RECT 222.85 36.47 224.73 36.63 ;
      RECT 224.57 35.86 224.73 36.63 ;
      RECT 223.71 35.23 223.87 36.63 ;
      RECT 222.85 35.86 223.01 36.63 ;
      RECT 224.67 35.23 224.83 36.05 ;
      RECT 222.75 35.23 222.91 36.05 ;
      RECT 224.67 37.11 224.83 38.19 ;
      RECT 223.71 36.79 223.87 38.19 ;
      RECT 222.75 37.11 222.91 38.19 ;
      RECT 224.57 36.79 224.73 37.39 ;
      RECT 222.85 36.79 223.01 37.39 ;
      RECT 222.85 36.79 224.73 36.95 ;
      RECT 223.47 50.66 223.63 51.5 ;
      RECT 223.47 50.66 224.27 50.82 ;
      RECT 224.11 50.18 224.27 50.82 ;
      RECT 224.11 50.18 224.75 50.5 ;
      RECT 224.59 47.07 224.75 50.5 ;
      RECT 224.27 47.07 224.75 47.23 ;
      RECT 224.27 45.44 224.43 47.23 ;
      RECT 224.59 56.67 224.75 61.86 ;
      RECT 223.31 56.67 224.75 56.83 ;
      RECT 224.43 54.4 224.59 56.83 ;
      RECT 223.31 56 223.47 56.83 ;
      RECT 224.27 47.39 224.43 49.72 ;
      RECT 223.95 47.39 224.43 47.55 ;
      RECT 223.95 43.85 224.11 47.55 ;
      RECT 223.95 43.85 224.73 44.01 ;
      RECT 224.57 39.56 224.73 44.01 ;
      RECT 224.39 39.56 224.73 39.84 ;
      RECT 224.39 39.16 224.55 39.84 ;
      RECT 223.17 53.23 223.45 53.51 ;
      RECT 223.29 53.03 223.45 53.51 ;
      RECT 223.29 53.03 224.27 53.19 ;
      RECT 224.11 50.98 224.27 53.19 ;
      RECT 224.11 52.54 224.31 52.82 ;
      RECT 224.11 50.98 224.65 51.14 ;
      RECT 224.43 50.8 224.65 51.14 ;
      RECT 222.83 68.07 224.65 68.23 ;
      RECT 224.49 62.02 224.65 68.23 ;
      RECT 224.27 62.02 224.65 62.18 ;
      RECT 224.27 57.45 224.43 62.18 ;
      RECT 222.83 57.45 224.43 57.61 ;
      RECT 222.83 57.39 223.15 57.61 ;
      RECT 222.99 53.74 223.15 57.61 ;
      RECT 222.83 51.32 222.99 53.9 ;
      RECT 222.83 51.32 223.31 51.48 ;
      RECT 223.15 49.88 223.31 51.48 ;
      RECT 223.15 49.88 223.63 50.04 ;
      RECT 223.47 47.71 223.63 50.04 ;
      RECT 223.47 47.71 224.09 47.99 ;
      RECT 224.11 54.06 224.27 56.51 ;
      RECT 224.11 54.06 224.63 54.22 ;
      RECT 224.47 51.34 224.63 54.22 ;
      RECT 224.43 52.98 224.63 54.22 ;
      RECT 224.43 51.34 224.63 52.12 ;
      RECT 224.07 34.44 224.41 34.72 ;
      RECT 224.07 32.44 224.23 34.72 ;
      RECT 224.07 33.11 224.41 33.39 ;
      RECT 224.07 32.44 224.41 32.72 ;
      RECT 224.07 40.7 224.41 40.98 ;
      RECT 224.07 38.7 224.23 40.98 ;
      RECT 224.07 40.03 224.41 40.31 ;
      RECT 224.07 38.7 224.41 38.98 ;
      RECT 223.71 55.68 223.87 56.51 ;
      RECT 223.47 55.68 223.87 55.84 ;
      RECT 223.47 53.67 223.63 55.84 ;
      RECT 223.47 53.67 224.11 53.83 ;
      RECT 223.83 53.35 224.11 53.83 ;
      RECT 223.57 51.7 223.95 51.92 ;
      RECT 223.79 50.98 223.95 51.92 ;
      RECT 223.15 52.58 223.91 52.86 ;
      RECT 223.75 52.18 223.91 52.86 ;
      RECT 223.15 51.64 223.31 52.86 ;
      RECT 223.47 62.9 223.63 67.89 ;
      RECT 223.47 65.82 223.69 66.55 ;
      RECT 223.15 47.39 223.31 49.72 ;
      RECT 223.15 47.39 223.63 47.55 ;
      RECT 223.47 43.85 223.63 47.55 ;
      RECT 222.85 43.85 223.63 44.01 ;
      RECT 222.85 39.56 223.01 44.01 ;
      RECT 222.85 39.56 223.19 39.84 ;
      RECT 223.03 39.16 223.19 39.84 ;
      RECT 223.17 34.44 223.51 34.72 ;
      RECT 223.35 32.44 223.51 34.72 ;
      RECT 223.17 33.11 223.51 33.39 ;
      RECT 223.17 32.44 223.51 32.72 ;
      RECT 223.17 40.7 223.51 40.98 ;
      RECT 223.35 38.7 223.51 40.98 ;
      RECT 223.17 40.03 223.51 40.31 ;
      RECT 223.17 38.7 223.51 38.98 ;
      RECT 222.99 62.9 223.15 67.89 ;
      RECT 222.99 64.59 223.27 65.31 ;
      RECT 222.51 46.75 222.67 47.43 ;
      RECT 222.19 46.75 222.99 46.91 ;
      RECT 222.83 44.23 222.99 46.91 ;
      RECT 222.19 44.23 222.35 46.91 ;
      RECT 221.99 10.08 222.15 11.89 ;
      RECT 221.99 10.08 222.73 10.24 ;
      RECT 222.51 8.88 222.67 10.24 ;
      RECT 222.51 7.5 222.67 8.72 ;
      RECT 222.46 7.58 222.67 7.9 ;
      RECT 221.43 7.59 222.67 7.75 ;
      RECT 222.39 7.58 222.67 7.75 ;
      RECT 214.47 15.8 214.63 16.08 ;
      RECT 211.35 15.8 211.51 16.08 ;
      RECT 213.87 15.8 214.63 15.96 ;
      RECT 211.35 15.8 212.11 15.96 ;
      RECT 211.95 14.07 212.11 15.96 ;
      RECT 220.37 14.25 220.53 15.89 ;
      RECT 205.45 14.25 205.61 15.89 ;
      RECT 212.91 12.21 213.07 15.8 ;
      RECT 213.87 14.07 214.03 15.96 ;
      RECT 217.85 14.12 218.03 15.79 ;
      RECT 216.57 14.1 216.73 15.79 ;
      RECT 209.25 14.1 209.41 15.79 ;
      RECT 207.95 14.12 208.13 15.79 ;
      RECT 221.71 14.64 221.87 15.6 ;
      RECT 204.11 14.64 204.27 15.6 ;
      RECT 222.51 12.64 222.67 14.96 ;
      RECT 203.31 12.64 203.47 14.96 ;
      RECT 215.53 14.1 215.69 14.89 ;
      RECT 210.29 14.1 210.45 14.89 ;
      RECT 220.09 14.64 222.67 14.84 ;
      RECT 203.31 14.64 205.89 14.84 ;
      RECT 205.73 12.56 205.89 14.84 ;
      RECT 220.09 14.25 221.54 14.84 ;
      RECT 204.44 14.25 205.89 14.84 ;
      RECT 214.59 14.36 215.69 14.52 ;
      RECT 210.29 14.36 211.39 14.52 ;
      RECT 211.23 14.08 211.39 14.52 ;
      RECT 214.59 14.08 214.75 14.52 ;
      RECT 216.57 14.12 220.25 14.28 ;
      RECT 204.44 14.25 209.41 14.28 ;
      RECT 215.53 14.1 217.05 14.26 ;
      RECT 208.93 14.1 210.45 14.26 ;
      RECT 205.73 14.12 210.45 14.26 ;
      RECT 213.87 14.08 214.75 14.24 ;
      RECT 211.23 14.08 212.11 14.24 ;
      RECT 211.77 14.07 214.21 14.23 ;
      RECT 220.09 12.56 220.25 14.84 ;
      RECT 219.13 12.55 219.29 14.28 ;
      RECT 218.25 13.45 218.41 14.28 ;
      RECT 207.57 13.45 207.73 14.28 ;
      RECT 206.69 12.55 206.85 14.28 ;
      RECT 215.79 12.32 215.95 14.26 ;
      RECT 210.03 12.32 210.19 14.26 ;
      RECT 214.05 13.38 214.21 14.24 ;
      RECT 211.77 13.38 211.93 14.24 ;
      RECT 218.17 12.55 218.33 13.61 ;
      RECT 207.65 12.55 207.81 13.61 ;
      RECT 213.93 13.38 214.21 13.54 ;
      RECT 211.77 13.38 212.05 13.54 ;
      RECT 221.84 17.18 222 18.9 ;
      RECT 221.84 17.96 222.67 18.12 ;
      RECT 222.51 17.84 222.67 18.12 ;
      RECT 221.8 17.06 221.96 17.34 ;
      RECT 220.82 19.61 220.98 21.25 ;
      RECT 213.87 20.42 214.03 21.25 ;
      RECT 212.91 16.39 213.07 21.25 ;
      RECT 211.95 20.42 212.11 21.25 ;
      RECT 205 19.61 205.16 21.25 ;
      RECT 221.6 20.89 222.02 21.05 ;
      RECT 219.86 19.61 220.02 21.05 ;
      RECT 205.96 19.61 206.12 21.05 ;
      RECT 203.96 20.89 204.38 21.05 ;
      RECT 204.22 19.61 204.38 21.05 ;
      RECT 218.86 20.21 219.02 20.89 ;
      RECT 216.61 20.43 216.77 20.89 ;
      RECT 209.21 20.43 209.37 20.89 ;
      RECT 206.96 20.21 207.12 20.89 ;
      RECT 221.6 19.61 221.76 21.05 ;
      RECT 216.15 20.43 216.77 20.59 ;
      RECT 209.21 20.43 209.83 20.59 ;
      RECT 209.67 19.1 209.83 20.59 ;
      RECT 213.95 19.16 214.11 20.58 ;
      RECT 211.87 19.16 212.03 20.58 ;
      RECT 215.19 19.16 215.35 20.49 ;
      RECT 210.63 19.16 210.79 20.49 ;
      RECT 216.15 19.1 216.31 20.59 ;
      RECT 218.86 20.21 220.02 20.37 ;
      RECT 219.82 19.61 220.02 20.37 ;
      RECT 205.96 20.21 207.12 20.37 ;
      RECT 205.96 19.61 206.16 20.37 ;
      RECT 219.82 19.61 220.98 19.81 ;
      RECT 205 19.61 206.16 19.81 ;
      RECT 219.65 19.61 222.59 19.77 ;
      RECT 203.39 19.61 206.33 19.77 ;
      RECT 206.17 19.1 206.33 19.77 ;
      RECT 218.69 19.1 218.97 19.73 ;
      RECT 207.01 19.1 207.29 19.73 ;
      RECT 219.65 19.1 219.81 19.77 ;
      RECT 215.19 19.16 216.31 19.37 ;
      RECT 209.67 19.16 210.79 19.37 ;
      RECT 209.67 19.16 216.31 19.32 ;
      RECT 215.3 19.1 219.81 19.26 ;
      RECT 214.83 18.46 214.99 19.32 ;
      RECT 213.87 17.56 214.03 19.32 ;
      RECT 211.95 17.56 212.11 19.32 ;
      RECT 210.99 18.46 211.15 19.32 ;
      RECT 206.17 19.1 210.68 19.26 ;
      RECT 209.54 17.76 209.7 19.26 ;
      RECT 216.28 19.01 218.2 19.26 ;
      RECT 218.02 16.65 218.2 19.26 ;
      RECT 207.78 19.01 209.7 19.26 ;
      RECT 217.08 17.58 217.24 19.26 ;
      RECT 216.28 17.76 216.44 19.26 ;
      RECT 208.74 17.58 208.9 19.26 ;
      RECT 207.78 16.65 207.96 19.26 ;
      RECT 215.75 17.76 216.44 17.92 ;
      RECT 209.54 17.76 210.23 17.92 ;
      RECT 210.07 16.77 210.23 17.92 ;
      RECT 215.75 16.77 215.91 17.92 ;
      RECT 222.28 15.57 222.44 17.28 ;
      RECT 221.68 16.43 221.84 16.71 ;
      RECT 221.68 16.43 222.44 16.59 ;
      RECT 222.22 15.57 222.5 15.73 ;
      RECT 220.29 34.88 222.49 35.04 ;
      RECT 222.21 34.59 222.49 35.04 ;
      RECT 221.27 34.59 221.51 35.04 ;
      RECT 220.29 34.59 220.57 35.04 ;
      RECT 221.27 38.38 221.51 39.02 ;
      RECT 222.21 38.38 222.49 38.83 ;
      RECT 220.29 38.38 220.57 38.83 ;
      RECT 220.29 38.38 222.49 38.54 ;
      RECT 221.81 23.66 222.35 23.82 ;
      RECT 222.19 20.12 222.35 23.82 ;
      RECT 221.89 23.22 222.35 23.38 ;
      RECT 222.19 20.83 222.44 21.11 ;
      RECT 221.92 20.12 222.35 20.28 ;
      RECT 222.24 26.15 222.4 28.96 ;
      RECT 222.24 26.15 222.43 26.51 ;
      RECT 220.45 36.47 222.33 36.63 ;
      RECT 222.17 35.88 222.33 36.63 ;
      RECT 221.31 35.23 221.47 36.63 ;
      RECT 220.45 35.88 220.61 36.63 ;
      RECT 222.27 35.23 222.43 36.06 ;
      RECT 220.35 35.23 220.51 36.06 ;
      RECT 222.27 37.11 222.43 38.19 ;
      RECT 221.31 36.79 221.47 38.19 ;
      RECT 220.35 37.11 220.51 38.19 ;
      RECT 222.17 36.79 222.33 37.39 ;
      RECT 220.45 36.79 220.61 37.39 ;
      RECT 220.45 36.79 222.33 36.95 ;
      RECT 220.53 68.07 222.35 68.23 ;
      RECT 220.53 62.02 220.69 68.23 ;
      RECT 220.53 62.02 220.91 62.18 ;
      RECT 220.75 57.45 220.91 62.18 ;
      RECT 220.75 57.45 222.35 57.61 ;
      RECT 222.03 57.39 222.35 57.61 ;
      RECT 222.03 53.74 222.19 57.61 ;
      RECT 222.19 51.32 222.35 53.9 ;
      RECT 221.87 51.32 222.35 51.48 ;
      RECT 221.87 49.88 222.03 51.48 ;
      RECT 221.55 49.88 222.03 50.04 ;
      RECT 221.55 47.71 221.71 50.04 ;
      RECT 221.09 47.71 221.71 47.99 ;
      RECT 221.87 47.39 222.03 49.72 ;
      RECT 221.55 47.39 222.03 47.55 ;
      RECT 221.55 43.85 221.71 47.55 ;
      RECT 221.55 43.85 222.33 44.01 ;
      RECT 222.17 39.56 222.33 44.01 ;
      RECT 221.99 39.56 222.33 39.84 ;
      RECT 221.99 39.16 222.15 39.84 ;
      RECT 219.69 8.96 220.01 9.12 ;
      RECT 219.69 7.8 219.85 9.12 ;
      RECT 222.03 7.91 222.19 8.8 ;
      RECT 221.11 7.91 222.19 8.07 ;
      RECT 219.69 7.8 221.27 7.96 ;
      RECT 222.01 23.98 222.19 24.52 ;
      RECT 221.49 23.98 222.19 24.14 ;
      RECT 221.49 23.27 221.65 24.14 ;
      RECT 221.55 21.78 221.71 23.43 ;
      RECT 221.41 21.21 221.57 21.94 ;
      RECT 221.28 20.95 221.44 21.37 ;
      RECT 222.03 62.9 222.19 67.89 ;
      RECT 221.91 64.59 222.19 65.31 ;
      RECT 221.27 52.58 222.03 52.86 ;
      RECT 221.87 51.64 222.03 52.86 ;
      RECT 221.27 52.18 221.43 52.86 ;
      RECT 221.67 34.44 222.01 34.72 ;
      RECT 221.67 32.44 221.83 34.72 ;
      RECT 221.67 33.11 222.01 33.39 ;
      RECT 221.67 32.44 222.01 32.72 ;
      RECT 221.67 40.7 222.01 40.98 ;
      RECT 221.67 38.7 221.83 40.98 ;
      RECT 221.67 40.03 222.01 40.31 ;
      RECT 221.67 38.7 222.01 38.98 ;
      RECT 221.73 53.23 222.01 53.51 ;
      RECT 221.73 53.03 221.89 53.51 ;
      RECT 220.91 53.03 221.89 53.19 ;
      RECT 220.91 50.98 221.07 53.19 ;
      RECT 220.87 52.54 221.07 52.82 ;
      RECT 220.53 50.98 221.07 51.14 ;
      RECT 220.53 50.8 220.75 51.14 ;
      RECT 220.91 28.52 222 28.68 ;
      RECT 220.91 28.35 221.19 28.68 ;
      RECT 220.51 28.35 221.19 28.51 ;
      RECT 221.76 24.79 221.92 28.32 ;
      RECT 221.23 25.16 221.92 25.32 ;
      RECT 221.71 12.92 221.87 13.67 ;
      RECT 221.51 12.92 221.87 13.08 ;
      RECT 221.51 9.68 221.67 13.08 ;
      RECT 221.51 9.68 221.71 11.89 ;
      RECT 220.73 9.68 221.71 9.84 ;
      RECT 220.73 8.6 220.89 9.84 ;
      RECT 220.43 56.67 220.59 61.86 ;
      RECT 220.43 56.67 221.87 56.83 ;
      RECT 221.71 56 221.87 56.83 ;
      RECT 220.59 54.4 220.75 56.83 ;
      RECT 219.87 26.02 220.43 26.18 ;
      RECT 220.27 25.58 220.43 26.18 ;
      RECT 220.27 25.58 220.97 25.74 ;
      RECT 220.81 22.71 220.97 25.74 ;
      RECT 220.77 24 220.97 25.74 ;
      RECT 220.77 24.3 221.77 24.46 ;
      RECT 220.71 22.04 220.87 22.99 ;
      RECT 220.55 21.85 220.71 22.32 ;
      RECT 221.55 50.66 221.71 51.5 ;
      RECT 220.91 50.66 221.71 50.82 ;
      RECT 220.91 50.18 221.07 50.82 ;
      RECT 220.43 50.18 221.07 50.5 ;
      RECT 220.43 47.07 220.59 50.5 ;
      RECT 220.43 47.07 220.91 47.23 ;
      RECT 220.75 45.44 220.91 47.23 ;
      RECT 221.31 55.68 221.47 56.51 ;
      RECT 221.31 55.68 221.71 55.84 ;
      RECT 221.55 53.67 221.71 55.84 ;
      RECT 221.07 53.67 221.71 53.83 ;
      RECT 221.07 53.35 221.35 53.83 ;
      RECT 221.55 62.9 221.71 67.89 ;
      RECT 221.49 65.82 221.71 66.55 ;
      RECT 221.23 51.7 221.61 51.92 ;
      RECT 221.23 50.98 221.39 51.92 ;
      RECT 218.65 26.36 218.81 26.72 ;
      RECT 218.65 26.36 220.95 26.52 ;
      RECT 220.79 26.04 220.95 26.52 ;
      RECT 220.79 26.04 221.6 26.2 ;
      RECT 221.36 16.52 221.52 18.9 ;
      RECT 221.16 16.52 221.52 16.8 ;
      RECT 221.23 15.31 221.39 16.8 ;
      RECT 221.03 22.13 221.39 22.41 ;
      RECT 221.03 21.53 221.19 22.41 ;
      RECT 220.16 21.53 220.32 21.92 ;
      RECT 220.16 21.53 221.19 21.69 ;
      RECT 220.34 20.21 220.5 21.69 ;
      RECT 221.19 11.5 221.35 13.22 ;
      RECT 219.83 12.22 221.35 12.38 ;
      RECT 220.93 11.5 221.35 11.66 ;
      RECT 220.75 47.39 220.91 49.72 ;
      RECT 220.75 47.39 221.23 47.55 ;
      RECT 221.07 43.85 221.23 47.55 ;
      RECT 220.45 43.85 221.23 44.01 ;
      RECT 220.45 39.56 220.61 44.01 ;
      RECT 220.45 39.56 220.79 39.84 ;
      RECT 220.63 39.16 220.79 39.84 ;
      RECT 220.26 18.3 221.2 18.46 ;
      RECT 220.84 17.05 221.2 18.46 ;
      RECT 220.84 16.2 221 18.46 ;
      RECT 220.09 16.2 221.05 16.36 ;
      RECT 220.89 16.08 221.05 16.36 ;
      RECT 219.65 16.07 220.32 16.23 ;
      RECT 220.77 34.44 221.11 34.72 ;
      RECT 220.95 32.44 221.11 34.72 ;
      RECT 220.77 33.11 221.11 33.39 ;
      RECT 220.77 32.44 221.11 32.72 ;
      RECT 220.77 40.7 221.11 40.98 ;
      RECT 220.95 38.7 221.11 40.98 ;
      RECT 220.77 40.03 221.11 40.31 ;
      RECT 220.77 38.7 221.11 38.98 ;
      RECT 220.91 54.06 221.07 56.51 ;
      RECT 220.55 54.06 221.07 54.22 ;
      RECT 220.55 52.98 220.75 54.22 ;
      RECT 220.55 51.34 220.71 54.22 ;
      RECT 220.55 51.34 220.75 52.12 ;
      RECT 218.82 28.01 220.98 28.17 ;
      RECT 220.82 26.68 220.98 28.17 ;
      RECT 219.82 26.97 219.98 28.17 ;
      RECT 218.82 27.93 219.14 28.17 ;
      RECT 218.82 27.34 218.98 28.17 ;
      RECT 219.61 12.56 219.77 13.61 ;
      RECT 219.51 11.9 219.67 13.24 ;
      RECT 219.51 11.9 220.79 12.06 ;
      RECT 219.69 9.6 219.85 12.06 ;
      RECT 220.5 16.52 220.68 16.84 ;
      RECT 219.78 16.52 220.68 16.68 ;
      RECT 220.49 23.18 220.65 23.84 ;
      RECT 220.32 23.18 220.65 23.34 ;
      RECT 220.32 22.65 220.48 23.34 ;
      RECT 220.11 46.75 220.27 47.43 ;
      RECT 219.79 46.75 220.59 46.91 ;
      RECT 220.43 44.23 220.59 46.91 ;
      RECT 219.79 44.23 219.95 46.91 ;
      RECT 220.3 26.69 220.46 27.85 ;
      RECT 220.26 26.69 220.5 27.33 ;
      RECT 220.17 9.28 220.33 11.72 ;
      RECT 219.21 8.12 219.37 11.72 ;
      RECT 218.25 8.5 218.41 11.72 ;
      RECT 216.59 9.63 216.75 11.4 ;
      RECT 216.59 9.95 218.41 10.11 ;
      RECT 217.28 9.79 217.44 10.11 ;
      RECT 220.21 8.12 220.41 9.84 ;
      RECT 216.53 9.63 217.04 9.79 ;
      RECT 219.21 9.28 220.41 9.44 ;
      RECT 218.21 8.5 218.52 8.78 ;
      RECT 218.21 8.56 219.37 8.72 ;
      RECT 215.23 28.74 220.35 28.9 ;
      RECT 218.43 27.92 218.59 28.9 ;
      RECT 216.99 27.92 217.15 28.9 ;
      RECT 220.04 16.92 220.2 18.12 ;
      RECT 219.8 16.92 220.2 17.08 ;
      RECT 217.89 34.88 220.09 35.04 ;
      RECT 219.81 34.59 220.09 35.04 ;
      RECT 218.87 34.59 219.11 35.04 ;
      RECT 217.89 34.59 218.17 35.04 ;
      RECT 218.87 38.38 219.11 39.02 ;
      RECT 219.81 38.38 220.09 38.83 ;
      RECT 217.89 38.38 218.17 38.83 ;
      RECT 217.89 38.38 220.09 38.54 ;
      RECT 217.71 21.69 217.87 26.21 ;
      RECT 218.95 24.34 219.11 26.2 ;
      RECT 216.47 24.35 216.63 26.2 ;
      RECT 219.83 24.04 220.05 25.52 ;
      RECT 215.53 24.04 215.75 25.52 ;
      RECT 218.95 24.46 220.05 24.63 ;
      RECT 215.53 24.46 216.63 24.63 ;
      RECT 216.45 21.69 216.61 24.63 ;
      RECT 218.97 21.69 219.13 24.63 ;
      RECT 216.45 21.69 219.13 21.85 ;
      RECT 218.05 36.47 219.93 36.63 ;
      RECT 219.77 35.86 219.93 36.63 ;
      RECT 218.91 35.23 219.07 36.63 ;
      RECT 218.05 35.86 218.21 36.63 ;
      RECT 219.87 35.23 220.03 36.05 ;
      RECT 217.95 35.23 218.11 36.05 ;
      RECT 219.87 37.11 220.03 38.19 ;
      RECT 218.91 36.79 219.07 38.19 ;
      RECT 217.95 37.11 218.11 38.19 ;
      RECT 219.77 36.79 219.93 37.39 ;
      RECT 218.05 36.79 218.21 37.39 ;
      RECT 218.05 36.79 219.93 36.95 ;
      RECT 219.83 21.37 219.99 23.37 ;
      RECT 215.99 21.37 219.99 21.53 ;
      RECT 219.34 20.73 219.5 21.53 ;
      RECT 215.99 20.78 216.15 21.53 ;
      RECT 218.67 50.66 218.83 51.5 ;
      RECT 218.67 50.66 219.47 50.82 ;
      RECT 219.31 50.18 219.47 50.82 ;
      RECT 219.31 50.18 219.95 50.5 ;
      RECT 219.79 47.07 219.95 50.5 ;
      RECT 219.47 47.07 219.95 47.23 ;
      RECT 219.47 45.44 219.63 47.23 ;
      RECT 219.79 56.67 219.95 61.86 ;
      RECT 218.51 56.67 219.95 56.83 ;
      RECT 219.63 54.4 219.79 56.83 ;
      RECT 218.51 56 218.67 56.83 ;
      RECT 219.47 47.39 219.63 49.72 ;
      RECT 219.15 47.39 219.63 47.55 ;
      RECT 219.15 43.85 219.31 47.55 ;
      RECT 219.15 43.85 219.93 44.01 ;
      RECT 219.77 39.56 219.93 44.01 ;
      RECT 219.59 39.56 219.93 39.84 ;
      RECT 219.59 39.16 219.75 39.84 ;
      RECT 218.37 53.23 218.65 53.51 ;
      RECT 218.49 53.03 218.65 53.51 ;
      RECT 218.49 53.03 219.47 53.19 ;
      RECT 219.31 50.98 219.47 53.19 ;
      RECT 219.31 52.54 219.51 52.82 ;
      RECT 219.31 50.98 219.85 51.14 ;
      RECT 219.63 50.8 219.85 51.14 ;
      RECT 218.03 68.07 219.85 68.23 ;
      RECT 219.69 62.02 219.85 68.23 ;
      RECT 219.47 62.02 219.85 62.18 ;
      RECT 219.47 57.45 219.63 62.18 ;
      RECT 218.03 57.45 219.63 57.61 ;
      RECT 218.03 57.39 218.35 57.61 ;
      RECT 218.19 53.74 218.35 57.61 ;
      RECT 218.03 51.32 218.19 53.9 ;
      RECT 218.03 51.32 218.51 51.48 ;
      RECT 218.35 49.88 218.51 51.48 ;
      RECT 218.35 49.88 218.83 50.04 ;
      RECT 218.67 47.71 218.83 50.04 ;
      RECT 218.67 47.71 219.29 47.99 ;
      RECT 219.31 54.06 219.47 56.51 ;
      RECT 219.31 54.06 219.83 54.22 ;
      RECT 219.67 51.34 219.83 54.22 ;
      RECT 219.63 52.98 219.83 54.22 ;
      RECT 219.63 51.34 219.83 52.12 ;
      RECT 218.52 18.78 219.64 18.94 ;
      RECT 219.46 17.48 219.64 18.94 ;
      RECT 217.56 17.26 217.73 18.8 ;
      RECT 217.57 16.12 217.73 18.8 ;
      RECT 216.6 16.44 216.76 18.8 ;
      RECT 218.52 16.03 218.68 18.94 ;
      RECT 216.55 16.44 216.76 17.57 ;
      RECT 219.46 16.44 219.62 18.94 ;
      RECT 216.55 17.26 217.73 17.42 ;
      RECT 216.55 16.44 216.83 17.42 ;
      RECT 219.33 14.52 219.49 16.71 ;
      RECT 215.55 16.12 218.68 16.28 ;
      RECT 218.37 14.52 218.53 16.28 ;
      RECT 217.37 14.84 217.53 16.28 ;
      RECT 218.37 14.52 219.49 14.68 ;
      RECT 219.27 34.44 219.61 34.72 ;
      RECT 219.27 32.44 219.43 34.72 ;
      RECT 219.27 33.11 219.61 33.39 ;
      RECT 219.27 32.44 219.61 32.72 ;
      RECT 219.27 40.7 219.61 40.98 ;
      RECT 219.27 38.7 219.43 40.98 ;
      RECT 219.27 40.03 219.61 40.31 ;
      RECT 219.27 38.7 219.61 38.98 ;
      RECT 219.43 21.85 219.59 24.3 ;
      RECT 219.29 21.85 219.59 22.13 ;
      RECT 219.27 24.79 219.47 25.35 ;
      RECT 219.27 24.79 219.59 25.03 ;
      RECT 217.95 28.04 218.27 28.32 ;
      RECT 218.11 25.99 218.27 28.32 ;
      RECT 219.3 27.02 219.46 27.7 ;
      RECT 218.11 27.02 219.46 27.18 ;
      RECT 218.11 25.99 218.49 26.23 ;
      RECT 218.33 25.16 218.49 26.23 ;
      RECT 217.97 20.26 218.13 21.05 ;
      RECT 217.97 20.26 218.7 20.44 ;
      RECT 218.54 19.89 218.7 20.44 ;
      RECT 218.54 19.89 219.36 20.05 ;
      RECT 219.17 19.61 219.36 20.05 ;
      RECT 219.17 19.61 219.45 19.77 ;
      RECT 218.91 55.68 219.07 56.51 ;
      RECT 218.67 55.68 219.07 55.84 ;
      RECT 218.67 53.67 218.83 55.84 ;
      RECT 218.67 53.67 219.31 53.83 ;
      RECT 219.03 53.35 219.31 53.83 ;
      RECT 218.77 51.7 219.15 51.92 ;
      RECT 218.99 50.98 219.15 51.92 ;
      RECT 218.35 52.58 219.11 52.86 ;
      RECT 218.95 52.18 219.11 52.86 ;
      RECT 218.35 51.64 218.51 52.86 ;
      RECT 218.65 12.53 218.81 13.61 ;
      RECT 218.81 11.88 218.97 12.69 ;
      RECT 217.85 11.77 218.09 12.05 ;
      RECT 217.85 11.88 218.97 12.04 ;
      RECT 218.73 8.88 218.89 12.04 ;
      RECT 218.67 62.9 218.83 67.89 ;
      RECT 218.67 65.82 218.89 66.55 ;
      RECT 218.35 47.39 218.51 49.72 ;
      RECT 218.35 47.39 218.83 47.55 ;
      RECT 218.67 43.85 218.83 47.55 ;
      RECT 218.05 43.85 218.83 44.01 ;
      RECT 218.05 39.56 218.21 44.01 ;
      RECT 218.05 39.56 218.39 39.84 ;
      RECT 218.23 39.16 218.39 39.84 ;
      RECT 218.65 22.01 218.81 23.37 ;
      RECT 218.03 22.01 218.81 22.17 ;
      RECT 218.33 24.72 218.71 24.96 ;
      RECT 218.33 22.35 218.49 24.96 ;
      RECT 218.37 34.44 218.71 34.72 ;
      RECT 218.55 32.44 218.71 34.72 ;
      RECT 218.37 33.11 218.71 33.39 ;
      RECT 218.37 32.44 218.71 32.72 ;
      RECT 218.37 40.7 218.71 40.98 ;
      RECT 218.55 38.7 218.71 40.98 ;
      RECT 218.37 40.03 218.71 40.31 ;
      RECT 218.37 38.7 218.71 38.98 ;
      RECT 217.07 12.21 217.23 13.28 ;
      RECT 217.07 12.21 218.65 12.37 ;
      RECT 217.53 11.47 217.69 12.37 ;
      RECT 217.59 10.85 217.75 11.63 ;
      RECT 218.19 62.9 218.35 67.89 ;
      RECT 218.19 64.59 218.47 65.31 ;
      RECT 217.71 46.75 217.87 47.43 ;
      RECT 217.39 46.75 218.19 46.91 ;
      RECT 218.03 44.23 218.19 46.91 ;
      RECT 217.39 44.23 217.55 46.91 ;
      RECT 217.91 10.51 218.07 11.24 ;
      RECT 217.41 10.51 218.07 10.67 ;
      RECT 217.76 8.96 217.92 9.79 ;
      RECT 216.73 8.96 217.92 9.12 ;
      RECT 217.43 20.63 217.71 20.79 ;
      RECT 217.55 19.59 217.71 20.79 ;
      RECT 215.49 34.88 217.69 35.04 ;
      RECT 217.41 34.59 217.69 35.04 ;
      RECT 216.47 34.59 216.71 35.04 ;
      RECT 215.49 34.59 215.77 35.04 ;
      RECT 216.47 38.38 216.71 39.02 ;
      RECT 217.41 38.38 217.69 38.83 ;
      RECT 215.49 38.38 215.77 38.83 ;
      RECT 215.49 38.38 217.69 38.54 ;
      RECT 217.31 28.04 217.63 28.32 ;
      RECT 217.31 25.99 217.47 28.32 ;
      RECT 216.12 27.02 216.28 27.7 ;
      RECT 216.12 27.02 217.47 27.18 ;
      RECT 217.09 25.99 217.47 26.23 ;
      RECT 217.09 25.16 217.25 26.23 ;
      RECT 215.65 36.47 217.53 36.63 ;
      RECT 217.37 35.88 217.53 36.63 ;
      RECT 216.51 35.23 216.67 36.63 ;
      RECT 215.65 35.88 215.81 36.63 ;
      RECT 217.47 35.23 217.63 36.06 ;
      RECT 215.55 35.23 215.71 36.06 ;
      RECT 217.47 37.11 217.63 38.19 ;
      RECT 216.51 36.79 216.67 38.19 ;
      RECT 215.55 37.11 215.71 38.19 ;
      RECT 217.37 36.79 217.53 37.39 ;
      RECT 215.65 36.79 215.81 37.39 ;
      RECT 215.65 36.79 217.53 36.95 ;
      RECT 216.77 22.01 216.93 23.37 ;
      RECT 216.77 22.01 217.55 22.17 ;
      RECT 215.73 68.07 217.55 68.23 ;
      RECT 215.73 62.02 215.89 68.23 ;
      RECT 215.73 62.02 216.11 62.18 ;
      RECT 215.95 57.45 216.11 62.18 ;
      RECT 215.95 57.45 217.55 57.61 ;
      RECT 217.23 57.39 217.55 57.61 ;
      RECT 217.23 53.74 217.39 57.61 ;
      RECT 217.39 51.32 217.55 53.9 ;
      RECT 217.07 51.32 217.55 51.48 ;
      RECT 217.07 49.88 217.23 51.48 ;
      RECT 216.75 49.88 217.23 50.04 ;
      RECT 216.75 47.71 216.91 50.04 ;
      RECT 216.29 47.71 216.91 47.99 ;
      RECT 217.07 47.39 217.23 49.72 ;
      RECT 216.75 47.39 217.23 47.55 ;
      RECT 216.75 43.85 216.91 47.55 ;
      RECT 216.75 43.85 217.53 44.01 ;
      RECT 217.37 39.56 217.53 44.01 ;
      RECT 217.19 39.56 217.53 39.84 ;
      RECT 217.19 39.16 217.35 39.84 ;
      RECT 216.89 14.44 217.05 15.64 ;
      RECT 216.89 14.44 217.39 14.6 ;
      RECT 217.23 62.9 217.39 67.89 ;
      RECT 217.11 64.59 217.39 65.31 ;
      RECT 216.87 24.72 217.25 24.96 ;
      RECT 217.09 22.35 217.25 24.96 ;
      RECT 216.59 12.32 216.75 13.37 ;
      RECT 216.71 11.56 216.87 12.48 ;
      RECT 216.11 11.56 217.23 11.72 ;
      RECT 217.07 10.27 217.23 11.72 ;
      RECT 216.11 10.4 216.27 11.72 ;
      RECT 216.47 52.58 217.23 52.86 ;
      RECT 217.07 51.64 217.23 52.86 ;
      RECT 216.47 52.18 216.63 52.86 ;
      RECT 216.87 34.44 217.21 34.72 ;
      RECT 216.87 32.44 217.03 34.72 ;
      RECT 216.87 33.11 217.21 33.39 ;
      RECT 216.87 32.44 217.21 32.72 ;
      RECT 216.87 40.7 217.21 40.98 ;
      RECT 216.87 38.7 217.03 40.98 ;
      RECT 216.87 40.03 217.21 40.31 ;
      RECT 216.87 38.7 217.21 38.98 ;
      RECT 216.93 53.23 217.21 53.51 ;
      RECT 216.93 53.03 217.09 53.51 ;
      RECT 216.11 53.03 217.09 53.19 ;
      RECT 216.11 50.98 216.27 53.19 ;
      RECT 216.07 52.54 216.27 52.82 ;
      RECT 215.73 50.98 216.27 51.14 ;
      RECT 215.73 50.8 215.95 51.14 ;
      RECT 215.63 56.67 215.79 61.86 ;
      RECT 215.63 56.67 217.07 56.83 ;
      RECT 216.91 56 217.07 56.83 ;
      RECT 215.79 54.4 215.95 56.83 ;
      RECT 216.77 26.36 216.93 26.72 ;
      RECT 214.63 26.36 216.93 26.52 ;
      RECT 214.63 26.04 214.79 26.52 ;
      RECT 213.98 26.04 214.79 26.2 ;
      RECT 216.75 50.66 216.91 51.5 ;
      RECT 216.11 50.66 216.91 50.82 ;
      RECT 216.11 50.18 216.27 50.82 ;
      RECT 215.63 50.18 216.27 50.5 ;
      RECT 215.63 47.07 215.79 50.5 ;
      RECT 215.63 47.07 216.11 47.23 ;
      RECT 215.95 45.44 216.11 47.23 ;
      RECT 216.51 55.68 216.67 56.51 ;
      RECT 216.51 55.68 216.91 55.84 ;
      RECT 216.75 53.67 216.91 55.84 ;
      RECT 216.27 53.67 216.91 53.83 ;
      RECT 216.27 53.35 216.55 53.83 ;
      RECT 216.75 62.9 216.91 67.89 ;
      RECT 216.69 65.82 216.91 66.55 ;
      RECT 216.43 51.7 216.81 51.92 ;
      RECT 216.43 50.98 216.59 51.92 ;
      RECT 214.6 28.01 216.76 28.17 ;
      RECT 216.6 27.34 216.76 28.17 ;
      RECT 216.44 27.93 216.76 28.17 ;
      RECT 215.6 26.97 215.76 28.17 ;
      RECT 214.6 26.68 214.76 28.17 ;
      RECT 216.11 12 216.27 12.84 ;
      RECT 216.11 12 216.55 12.16 ;
      RECT 216.39 11.88 216.55 12.16 ;
      RECT 214.86 8.82 216.45 8.98 ;
      RECT 216.29 7.16 216.45 8.98 ;
      RECT 215.95 47.39 216.11 49.72 ;
      RECT 215.95 47.39 216.43 47.55 ;
      RECT 216.27 43.85 216.43 47.55 ;
      RECT 215.65 43.85 216.43 44.01 ;
      RECT 215.65 39.56 215.81 44.01 ;
      RECT 215.65 39.56 215.99 39.84 ;
      RECT 215.83 39.16 215.99 39.84 ;
      RECT 216.26 9.92 216.42 10.24 ;
      RECT 216.02 9.92 216.42 10.12 ;
      RECT 215.23 15.8 215.39 17.77 ;
      RECT 215.23 15.8 216.05 15.96 ;
      RECT 216.05 14.42 216.21 15.88 ;
      RECT 215.87 15.72 216.21 15.88 ;
      RECT 216.05 14.42 216.39 14.58 ;
      RECT 216.11 24.79 216.31 25.35 ;
      RECT 215.99 24.79 216.31 25.03 ;
      RECT 215.97 34.44 216.31 34.72 ;
      RECT 216.15 32.44 216.31 34.72 ;
      RECT 215.97 33.11 216.31 33.39 ;
      RECT 215.97 32.44 216.31 32.72 ;
      RECT 215.97 40.7 216.31 40.98 ;
      RECT 216.15 38.7 216.31 40.98 ;
      RECT 215.97 40.03 216.31 40.31 ;
      RECT 215.97 38.7 216.31 38.98 ;
      RECT 215.99 21.85 216.15 24.3 ;
      RECT 215.99 21.85 216.29 22.13 ;
      RECT 216.11 54.06 216.27 56.51 ;
      RECT 215.75 54.06 216.27 54.22 ;
      RECT 215.75 52.98 215.95 54.22 ;
      RECT 215.75 51.34 215.91 54.22 ;
      RECT 215.75 51.34 215.95 52.12 ;
      RECT 215.61 18.51 215.8 18.94 ;
      RECT 215.41 18.51 216.1 18.7 ;
      RECT 215.59 21.29 215.75 23.37 ;
      RECT 215.67 19.81 215.83 21.46 ;
      RECT 215.21 12.58 215.49 13.24 ;
      RECT 215.33 11.84 215.49 13.24 ;
      RECT 214.97 11.84 215.13 12.12 ;
      RECT 214.97 11.84 215.81 12 ;
      RECT 215.65 10.46 215.81 12 ;
      RECT 215.31 46.75 215.47 47.43 ;
      RECT 214.99 46.75 215.79 46.91 ;
      RECT 215.63 44.23 215.79 46.91 ;
      RECT 214.99 44.23 215.15 46.91 ;
      RECT 215.15 26.02 215.71 26.18 ;
      RECT 215.15 25.58 215.31 26.18 ;
      RECT 214.61 25.58 215.31 25.74 ;
      RECT 214.61 24 214.81 25.74 ;
      RECT 213.87 24.24 214.81 24.52 ;
      RECT 213.87 21.85 214.03 24.52 ;
      RECT 214.54 9.14 214.73 9.52 ;
      RECT 214.54 9.14 215.67 9.3 ;
      RECT 214.54 8.52 214.7 9.52 ;
      RECT 214.52 8.36 214.68 8.64 ;
      RECT 214.91 18.13 215.57 18.3 ;
      RECT 214.91 15 215.07 18.3 ;
      RECT 214.91 15.32 215.61 15.64 ;
      RECT 214.45 15 215.07 15.16 ;
      RECT 215.17 9.68 215.33 11.68 ;
      RECT 210.65 9.68 210.81 11.68 ;
      RECT 213.71 9.68 213.87 11.36 ;
      RECT 212.11 9.68 212.27 11.36 ;
      RECT 212.11 10.76 213.87 10.92 ;
      RECT 212.91 8.38 213.07 10.92 ;
      RECT 213.71 9.68 215.33 9.84 ;
      RECT 215.05 9.46 215.21 9.84 ;
      RECT 210.65 9.68 212.27 9.84 ;
      RECT 210.77 9.46 210.93 9.84 ;
      RECT 215.12 26.68 215.28 27.85 ;
      RECT 215.08 26.68 215.32 27.33 ;
      RECT 213.09 34.88 215.29 35.04 ;
      RECT 215.01 34.59 215.29 35.04 ;
      RECT 214.07 34.59 214.31 35.04 ;
      RECT 213.09 34.59 213.37 35.04 ;
      RECT 214.07 38.38 214.31 39.02 ;
      RECT 215.01 38.38 215.29 38.83 ;
      RECT 213.09 38.38 213.37 38.83 ;
      RECT 213.09 38.38 215.29 38.54 ;
      RECT 215.07 13.5 215.23 14.2 ;
      RECT 214.89 13.5 215.23 13.66 ;
      RECT 214.89 12.52 215.05 13.66 ;
      RECT 214.65 12.52 215.05 12.84 ;
      RECT 214.65 10.84 214.81 12.84 ;
      RECT 213.25 36.47 215.13 36.63 ;
      RECT 214.97 35.86 215.13 36.63 ;
      RECT 214.11 35.23 214.27 36.63 ;
      RECT 213.25 35.86 213.41 36.63 ;
      RECT 215.07 35.23 215.23 36.05 ;
      RECT 213.15 35.23 213.31 36.05 ;
      RECT 215.07 37.11 215.23 38.19 ;
      RECT 214.11 36.79 214.27 38.19 ;
      RECT 213.15 37.11 213.31 38.19 ;
      RECT 214.97 36.79 215.13 37.39 ;
      RECT 213.25 36.79 213.41 37.39 ;
      RECT 213.25 36.79 215.13 36.95 ;
      RECT 213.87 50.66 214.03 51.5 ;
      RECT 213.87 50.66 214.67 50.82 ;
      RECT 214.51 50.18 214.67 50.82 ;
      RECT 214.51 50.18 215.15 50.5 ;
      RECT 214.99 47.07 215.15 50.5 ;
      RECT 214.67 47.07 215.15 47.23 ;
      RECT 214.67 45.44 214.83 47.23 ;
      RECT 214.99 56.67 215.15 61.86 ;
      RECT 213.71 56.67 215.15 56.83 ;
      RECT 214.83 54.4 214.99 56.83 ;
      RECT 213.71 56 213.87 56.83 ;
      RECT 214.67 47.39 214.83 49.72 ;
      RECT 214.35 47.39 214.83 47.55 ;
      RECT 214.35 43.85 214.51 47.55 ;
      RECT 214.35 43.85 215.13 44.01 ;
      RECT 214.97 39.56 215.13 44.01 ;
      RECT 214.79 39.56 215.13 39.84 ;
      RECT 214.79 39.16 214.95 39.84 ;
      RECT 214.93 23.12 215.09 23.84 ;
      RECT 214.19 23.12 215.09 23.28 ;
      RECT 214.19 20.86 214.35 23.28 ;
      RECT 214.19 20.86 214.55 21.02 ;
      RECT 214.39 20.74 214.55 21.02 ;
      RECT 213.58 28.52 214.67 28.68 ;
      RECT 214.39 28.35 214.67 28.68 ;
      RECT 214.39 28.35 215.07 28.51 ;
      RECT 213.57 53.23 213.85 53.51 ;
      RECT 213.69 53.03 213.85 53.51 ;
      RECT 213.69 53.03 214.67 53.19 ;
      RECT 214.51 50.98 214.67 53.19 ;
      RECT 214.51 52.54 214.71 52.82 ;
      RECT 214.51 50.98 215.05 51.14 ;
      RECT 214.83 50.8 215.05 51.14 ;
      RECT 213.23 68.07 215.05 68.23 ;
      RECT 214.89 62.02 215.05 68.23 ;
      RECT 214.67 62.02 215.05 62.18 ;
      RECT 214.67 57.45 214.83 62.18 ;
      RECT 213.23 57.45 214.83 57.61 ;
      RECT 213.23 57.39 213.55 57.61 ;
      RECT 213.39 53.74 213.55 57.61 ;
      RECT 213.23 51.32 213.39 53.9 ;
      RECT 213.23 51.32 213.71 51.48 ;
      RECT 213.55 49.88 213.71 51.48 ;
      RECT 213.55 49.88 214.03 50.04 ;
      RECT 213.87 47.71 214.03 50.04 ;
      RECT 213.87 47.71 214.49 47.99 ;
      RECT 214.51 54.06 214.67 56.51 ;
      RECT 214.51 54.06 215.03 54.22 ;
      RECT 214.87 51.34 215.03 54.22 ;
      RECT 214.83 52.98 215.03 54.22 ;
      RECT 214.83 51.34 215.03 52.12 ;
      RECT 214.47 13.06 214.63 13.54 ;
      RECT 214.19 13.06 214.63 13.22 ;
      RECT 214.19 10 214.35 13.22 ;
      RECT 214.19 10 215.01 10.16 ;
      RECT 214.55 22.29 214.79 22.53 ;
      RECT 214.55 21.18 214.71 22.53 ;
      RECT 214.51 21.18 214.71 21.58 ;
      RECT 214.71 19.81 214.88 21.35 ;
      RECT 214.47 34.44 214.81 34.72 ;
      RECT 214.47 32.44 214.63 34.72 ;
      RECT 214.47 33.11 214.81 33.39 ;
      RECT 214.47 32.44 214.81 32.72 ;
      RECT 214.47 40.7 214.81 40.98 ;
      RECT 214.47 38.7 214.63 40.98 ;
      RECT 214.47 40.03 214.81 40.31 ;
      RECT 214.47 38.7 214.81 38.98 ;
      RECT 214.35 17.24 214.51 19 ;
      RECT 213.39 14.39 213.55 18.85 ;
      RECT 213.39 17.24 214.51 17.4 ;
      RECT 213.37 15.32 213.57 16.04 ;
      RECT 213.39 14.39 213.57 16.04 ;
      RECT 214.11 55.68 214.27 56.51 ;
      RECT 213.87 55.68 214.27 55.84 ;
      RECT 213.87 53.67 214.03 55.84 ;
      RECT 213.87 53.67 214.51 53.83 ;
      RECT 214.23 53.35 214.51 53.83 ;
      RECT 213.66 24.7 213.82 28.32 ;
      RECT 213.66 25.16 214.35 25.32 ;
      RECT 213.13 24.7 213.82 24.86 ;
      RECT 213.97 51.7 214.35 51.92 ;
      RECT 214.19 50.98 214.35 51.92 ;
      RECT 213.55 52.58 214.31 52.86 ;
      RECT 214.15 52.18 214.31 52.86 ;
      RECT 213.55 51.64 213.71 52.86 ;
      RECT 213.87 62.9 214.03 67.89 ;
      RECT 213.87 65.82 214.09 66.55 ;
      RECT 213.31 9.36 213.47 10.6 ;
      RECT 213.31 9.36 214.05 9.52 ;
      RECT 213.55 47.39 213.71 49.72 ;
      RECT 213.55 47.39 214.03 47.55 ;
      RECT 213.87 43.85 214.03 47.55 ;
      RECT 213.25 43.85 214.03 44.01 ;
      RECT 213.25 39.56 213.41 44.01 ;
      RECT 213.25 39.56 213.59 39.84 ;
      RECT 213.43 39.16 213.59 39.84 ;
      RECT 213.57 34.44 213.91 34.72 ;
      RECT 213.75 32.44 213.91 34.72 ;
      RECT 213.57 33.11 213.91 33.39 ;
      RECT 213.57 32.44 213.91 32.72 ;
      RECT 213.57 40.7 213.91 40.98 ;
      RECT 213.75 38.7 213.91 40.98 ;
      RECT 213.57 40.03 213.91 40.31 ;
      RECT 213.57 38.7 213.91 38.98 ;
      RECT 213.47 11.52 213.63 12.43 ;
      RECT 213.47 11.75 213.71 12.03 ;
      RECT 213.19 11.52 213.63 11.68 ;
      RECT 213.19 11.08 213.35 11.68 ;
      RECT 213.39 62.9 213.55 67.89 ;
      RECT 213.39 64.59 213.67 65.31 ;
      RECT 213.39 23.73 213.57 24.54 ;
      RECT 213.39 20.48 213.55 24.54 ;
      RECT 212.91 46.75 213.07 47.43 ;
      RECT 212.59 46.75 213.39 46.91 ;
      RECT 213.23 44.23 213.39 46.91 ;
      RECT 212.59 44.23 212.75 46.91 ;
      RECT 213.18 26.15 213.34 28.96 ;
      RECT 213.15 26.15 213.34 26.51 ;
      RECT 210.69 34.88 212.89 35.04 ;
      RECT 212.61 34.59 212.89 35.04 ;
      RECT 211.67 34.59 211.91 35.04 ;
      RECT 210.69 34.59 210.97 35.04 ;
      RECT 211.67 38.38 211.91 39.02 ;
      RECT 212.61 38.38 212.89 38.83 ;
      RECT 210.69 38.38 210.97 38.83 ;
      RECT 210.69 38.38 212.89 38.54 ;
      RECT 212.16 24.7 212.32 28.32 ;
      RECT 211.63 25.16 212.32 25.32 ;
      RECT 212.16 24.7 212.85 24.86 ;
      RECT 212.64 26.15 212.8 28.96 ;
      RECT 212.64 26.15 212.83 26.51 ;
      RECT 210.85 36.47 212.73 36.63 ;
      RECT 212.57 35.88 212.73 36.63 ;
      RECT 211.71 35.23 211.87 36.63 ;
      RECT 210.85 35.88 211.01 36.63 ;
      RECT 212.67 35.23 212.83 36.06 ;
      RECT 210.75 35.23 210.91 36.06 ;
      RECT 212.67 37.11 212.83 38.19 ;
      RECT 211.71 36.79 211.87 38.19 ;
      RECT 210.75 37.11 210.91 38.19 ;
      RECT 212.57 36.79 212.73 37.39 ;
      RECT 210.85 36.79 211.01 37.39 ;
      RECT 210.85 36.79 212.73 36.95 ;
      RECT 212.35 11.52 212.51 12.43 ;
      RECT 212.27 11.75 212.51 12.03 ;
      RECT 212.35 11.52 212.79 11.68 ;
      RECT 212.63 11.08 212.79 11.68 ;
      RECT 210.93 68.07 212.75 68.23 ;
      RECT 210.93 62.02 211.09 68.23 ;
      RECT 210.93 62.02 211.31 62.18 ;
      RECT 211.15 57.45 211.31 62.18 ;
      RECT 211.15 57.45 212.75 57.61 ;
      RECT 212.43 57.39 212.75 57.61 ;
      RECT 212.43 53.74 212.59 57.61 ;
      RECT 212.59 51.32 212.75 53.9 ;
      RECT 212.27 51.32 212.75 51.48 ;
      RECT 212.27 49.88 212.43 51.48 ;
      RECT 211.95 49.88 212.43 50.04 ;
      RECT 211.95 47.71 212.11 50.04 ;
      RECT 211.49 47.71 212.11 47.99 ;
      RECT 212.27 47.39 212.43 49.72 ;
      RECT 211.95 47.39 212.43 47.55 ;
      RECT 211.95 43.85 212.11 47.55 ;
      RECT 211.95 43.85 212.73 44.01 ;
      RECT 212.57 39.56 212.73 44.01 ;
      RECT 212.39 39.56 212.73 39.84 ;
      RECT 212.39 39.16 212.55 39.84 ;
      RECT 212.51 9.36 212.67 10.6 ;
      RECT 211.93 9.36 212.67 9.52 ;
      RECT 211.47 17.24 211.63 19 ;
      RECT 212.43 14.39 212.59 18.85 ;
      RECT 211.47 17.24 212.59 17.4 ;
      RECT 212.41 15.32 212.61 16.04 ;
      RECT 212.41 14.39 212.59 16.04 ;
      RECT 212.41 23.73 212.59 24.54 ;
      RECT 212.43 20.48 212.59 24.54 ;
      RECT 212.43 62.9 212.59 67.89 ;
      RECT 212.31 64.59 212.59 65.31 ;
      RECT 211.67 52.58 212.43 52.86 ;
      RECT 212.27 51.64 212.43 52.86 ;
      RECT 211.67 52.18 211.83 52.86 ;
      RECT 212.07 34.44 212.41 34.72 ;
      RECT 212.07 32.44 212.23 34.72 ;
      RECT 212.07 33.11 212.41 33.39 ;
      RECT 212.07 32.44 212.41 32.72 ;
      RECT 212.07 40.7 212.41 40.98 ;
      RECT 212.07 38.7 212.23 40.98 ;
      RECT 212.07 40.03 212.41 40.31 ;
      RECT 212.07 38.7 212.41 38.98 ;
      RECT 212.13 53.23 212.41 53.51 ;
      RECT 212.13 53.03 212.29 53.51 ;
      RECT 211.31 53.03 212.29 53.19 ;
      RECT 211.31 50.98 211.47 53.19 ;
      RECT 211.27 52.54 211.47 52.82 ;
      RECT 210.93 50.98 211.47 51.14 ;
      RECT 210.93 50.8 211.15 51.14 ;
      RECT 211.31 28.52 212.4 28.68 ;
      RECT 211.31 28.35 211.59 28.68 ;
      RECT 210.91 28.35 211.59 28.51 ;
      RECT 210.83 56.67 210.99 61.86 ;
      RECT 210.83 56.67 212.27 56.83 ;
      RECT 212.11 56 212.27 56.83 ;
      RECT 210.99 54.4 211.15 56.83 ;
      RECT 210.27 26.02 210.83 26.18 ;
      RECT 210.67 25.58 210.83 26.18 ;
      RECT 210.67 25.58 211.37 25.74 ;
      RECT 211.17 24 211.37 25.74 ;
      RECT 211.17 24.24 212.11 24.52 ;
      RECT 211.95 21.85 212.11 24.52 ;
      RECT 211.95 50.66 212.11 51.5 ;
      RECT 211.31 50.66 212.11 50.82 ;
      RECT 211.31 50.18 211.47 50.82 ;
      RECT 210.83 50.18 211.47 50.5 ;
      RECT 210.83 47.07 210.99 50.5 ;
      RECT 210.83 47.07 211.31 47.23 ;
      RECT 211.15 45.44 211.31 47.23 ;
      RECT 211.71 55.68 211.87 56.51 ;
      RECT 211.71 55.68 212.11 55.84 ;
      RECT 211.95 53.67 212.11 55.84 ;
      RECT 211.47 53.67 212.11 53.83 ;
      RECT 211.47 53.35 211.75 53.83 ;
      RECT 211.95 62.9 212.11 67.89 ;
      RECT 211.89 65.82 212.11 66.55 ;
      RECT 211.63 51.7 212.01 51.92 ;
      RECT 211.63 50.98 211.79 51.92 ;
      RECT 209.05 26.36 209.21 26.72 ;
      RECT 209.05 26.36 211.35 26.52 ;
      RECT 211.19 26.04 211.35 26.52 ;
      RECT 211.19 26.04 212 26.2 ;
      RECT 211.35 13.06 211.51 13.54 ;
      RECT 211.35 13.06 211.79 13.22 ;
      RECT 211.63 10 211.79 13.22 ;
      RECT 210.97 10 211.79 10.16 ;
      RECT 210.89 23.12 211.05 23.84 ;
      RECT 210.89 23.12 211.79 23.28 ;
      RECT 211.63 20.86 211.79 23.28 ;
      RECT 211.43 20.86 211.79 21.02 ;
      RECT 211.43 20.74 211.59 21.02 ;
      RECT 211.15 47.39 211.31 49.72 ;
      RECT 211.15 47.39 211.63 47.55 ;
      RECT 211.47 43.85 211.63 47.55 ;
      RECT 210.85 43.85 211.63 44.01 ;
      RECT 210.85 39.56 211.01 44.01 ;
      RECT 210.85 39.56 211.19 39.84 ;
      RECT 211.03 39.16 211.19 39.84 ;
      RECT 210.41 18.13 211.07 18.3 ;
      RECT 210.91 15 211.07 18.3 ;
      RECT 210.37 15.32 211.07 15.64 ;
      RECT 210.91 15 211.53 15.16 ;
      RECT 211.17 34.44 211.51 34.72 ;
      RECT 211.35 32.44 211.51 34.72 ;
      RECT 211.17 33.11 211.51 33.39 ;
      RECT 211.17 32.44 211.51 32.72 ;
      RECT 211.17 40.7 211.51 40.98 ;
      RECT 211.35 38.7 211.51 40.98 ;
      RECT 211.17 40.03 211.51 40.31 ;
      RECT 211.17 38.7 211.51 38.98 ;
      RECT 211.19 22.29 211.43 22.53 ;
      RECT 211.27 21.18 211.43 22.53 ;
      RECT 211.27 21.18 211.47 21.58 ;
      RECT 211.1 19.81 211.27 21.35 ;
      RECT 211.31 54.06 211.47 56.51 ;
      RECT 210.95 54.06 211.47 54.22 ;
      RECT 210.95 52.98 211.15 54.22 ;
      RECT 210.95 51.34 211.11 54.22 ;
      RECT 210.95 51.34 211.15 52.12 ;
      RECT 211.25 9.14 211.44 9.52 ;
      RECT 210.31 9.14 211.44 9.3 ;
      RECT 211.28 8.52 211.44 9.52 ;
      RECT 211.3 8.36 211.46 8.64 ;
      RECT 209.22 28.01 211.38 28.17 ;
      RECT 211.22 26.68 211.38 28.17 ;
      RECT 210.22 26.97 210.38 28.17 ;
      RECT 209.22 27.93 209.54 28.17 ;
      RECT 209.22 27.34 209.38 28.17 ;
      RECT 210.75 13.5 210.91 14.2 ;
      RECT 210.75 13.5 211.09 13.66 ;
      RECT 210.93 12.52 211.09 13.66 ;
      RECT 210.93 12.52 211.33 12.84 ;
      RECT 211.17 10.84 211.33 12.84 ;
      RECT 209.53 8.82 211.12 8.98 ;
      RECT 209.53 7.16 209.69 8.98 ;
      RECT 210.49 12.58 210.77 13.24 ;
      RECT 210.49 11.84 210.65 13.24 ;
      RECT 210.85 11.84 211.01 12.12 ;
      RECT 210.17 11.84 211.01 12 ;
      RECT 210.17 10.46 210.33 12 ;
      RECT 210.51 46.75 210.67 47.43 ;
      RECT 210.19 46.75 210.99 46.91 ;
      RECT 210.83 44.23 210.99 46.91 ;
      RECT 210.19 44.23 210.35 46.91 ;
      RECT 210.7 26.68 210.86 27.85 ;
      RECT 210.66 26.68 210.9 27.33 ;
      RECT 210.59 15.8 210.75 17.77 ;
      RECT 209.93 15.8 210.75 15.96 ;
      RECT 209.77 14.42 209.93 15.88 ;
      RECT 209.77 15.72 210.11 15.88 ;
      RECT 209.59 14.42 209.93 14.58 ;
      RECT 205.63 28.74 210.75 28.9 ;
      RECT 208.83 27.92 208.99 28.9 ;
      RECT 207.39 27.92 207.55 28.9 ;
      RECT 210.18 18.51 210.37 18.94 ;
      RECT 209.88 18.51 210.57 18.7 ;
      RECT 208.29 34.88 210.49 35.04 ;
      RECT 210.21 34.59 210.49 35.04 ;
      RECT 209.27 34.59 209.51 35.04 ;
      RECT 208.29 34.59 208.57 35.04 ;
      RECT 209.27 38.38 209.51 39.02 ;
      RECT 210.21 38.38 210.49 38.83 ;
      RECT 208.29 38.38 208.57 38.83 ;
      RECT 208.29 38.38 210.49 38.54 ;
      RECT 208.11 21.69 208.27 26.21 ;
      RECT 209.35 24.35 209.51 26.2 ;
      RECT 206.87 24.34 207.03 26.2 ;
      RECT 210.23 24.04 210.45 25.52 ;
      RECT 205.93 24.04 206.15 25.52 ;
      RECT 209.35 24.46 210.45 24.63 ;
      RECT 205.93 24.46 207.03 24.63 ;
      RECT 206.85 21.69 207.01 24.63 ;
      RECT 209.37 21.69 209.53 24.63 ;
      RECT 206.85 21.69 209.53 21.85 ;
      RECT 206.34 18.78 207.46 18.94 ;
      RECT 209.22 16.44 209.38 18.8 ;
      RECT 208.25 17.26 208.42 18.8 ;
      RECT 207.3 16.03 207.46 18.94 ;
      RECT 206.34 17.48 206.52 18.94 ;
      RECT 209.22 16.44 209.43 17.57 ;
      RECT 206.36 16.44 206.52 18.94 ;
      RECT 208.25 17.26 209.43 17.42 ;
      RECT 209.15 16.44 209.43 17.42 ;
      RECT 208.25 16.12 208.41 18.8 ;
      RECT 206.49 14.52 206.65 16.71 ;
      RECT 207.3 16.12 210.43 16.28 ;
      RECT 208.45 14.84 208.61 16.28 ;
      RECT 207.45 14.52 207.61 16.28 ;
      RECT 206.49 14.52 207.61 14.68 ;
      RECT 208.45 36.47 210.33 36.63 ;
      RECT 210.17 35.86 210.33 36.63 ;
      RECT 209.31 35.23 209.47 36.63 ;
      RECT 208.45 35.86 208.61 36.63 ;
      RECT 210.27 35.23 210.43 36.05 ;
      RECT 208.35 35.23 208.51 36.05 ;
      RECT 210.27 37.11 210.43 38.19 ;
      RECT 209.31 36.79 209.47 38.19 ;
      RECT 208.35 37.11 208.51 38.19 ;
      RECT 210.17 36.79 210.33 37.39 ;
      RECT 208.45 36.79 208.61 37.39 ;
      RECT 208.45 36.79 210.33 36.95 ;
      RECT 210.23 21.29 210.39 23.37 ;
      RECT 210.15 19.81 210.31 21.46 ;
      RECT 209.07 50.66 209.23 51.5 ;
      RECT 209.07 50.66 209.87 50.82 ;
      RECT 209.71 50.18 209.87 50.82 ;
      RECT 209.71 50.18 210.35 50.5 ;
      RECT 210.19 47.07 210.35 50.5 ;
      RECT 209.87 47.07 210.35 47.23 ;
      RECT 209.87 45.44 210.03 47.23 ;
      RECT 210.19 56.67 210.35 61.86 ;
      RECT 208.91 56.67 210.35 56.83 ;
      RECT 210.03 54.4 210.19 56.83 ;
      RECT 208.91 56 209.07 56.83 ;
      RECT 209.87 47.39 210.03 49.72 ;
      RECT 209.55 47.39 210.03 47.55 ;
      RECT 209.55 43.85 209.71 47.55 ;
      RECT 209.55 43.85 210.33 44.01 ;
      RECT 210.17 39.56 210.33 44.01 ;
      RECT 209.99 39.56 210.33 39.84 ;
      RECT 209.99 39.16 210.15 39.84 ;
      RECT 208.77 53.23 209.05 53.51 ;
      RECT 208.89 53.03 209.05 53.51 ;
      RECT 208.89 53.03 209.87 53.19 ;
      RECT 209.71 50.98 209.87 53.19 ;
      RECT 209.71 52.54 209.91 52.82 ;
      RECT 209.71 50.98 210.25 51.14 ;
      RECT 210.03 50.8 210.25 51.14 ;
      RECT 208.43 68.07 210.25 68.23 ;
      RECT 210.09 62.02 210.25 68.23 ;
      RECT 209.87 62.02 210.25 62.18 ;
      RECT 209.87 57.45 210.03 62.18 ;
      RECT 208.43 57.45 210.03 57.61 ;
      RECT 208.43 57.39 208.75 57.61 ;
      RECT 208.59 53.74 208.75 57.61 ;
      RECT 208.43 51.32 208.59 53.9 ;
      RECT 208.43 51.32 208.91 51.48 ;
      RECT 208.75 49.88 208.91 51.48 ;
      RECT 208.75 49.88 209.23 50.04 ;
      RECT 209.07 47.71 209.23 50.04 ;
      RECT 209.07 47.71 209.69 47.99 ;
      RECT 209.71 54.06 209.87 56.51 ;
      RECT 209.71 54.06 210.23 54.22 ;
      RECT 210.07 51.34 210.23 54.22 ;
      RECT 210.03 52.98 210.23 54.22 ;
      RECT 210.03 51.34 210.23 52.12 ;
      RECT 209.67 34.44 210.01 34.72 ;
      RECT 209.67 32.44 209.83 34.72 ;
      RECT 209.67 33.11 210.01 33.39 ;
      RECT 209.67 32.44 210.01 32.72 ;
      RECT 209.67 40.7 210.01 40.98 ;
      RECT 209.67 38.7 209.83 40.98 ;
      RECT 209.67 40.03 210.01 40.31 ;
      RECT 209.67 38.7 210.01 38.98 ;
      RECT 205.99 21.37 206.15 23.37 ;
      RECT 205.99 21.37 209.99 21.53 ;
      RECT 209.83 20.78 209.99 21.53 ;
      RECT 206.48 20.73 206.64 21.53 ;
      RECT 209.83 21.85 209.99 24.3 ;
      RECT 209.69 21.85 209.99 22.13 ;
      RECT 209.67 24.79 209.87 25.35 ;
      RECT 209.67 24.79 209.99 25.03 ;
      RECT 209.56 9.92 209.72 10.24 ;
      RECT 209.56 9.92 209.96 10.12 ;
      RECT 209.23 12.32 209.39 13.37 ;
      RECT 209.11 11.56 209.27 12.48 ;
      RECT 208.75 11.56 209.87 11.72 ;
      RECT 209.71 10.4 209.87 11.72 ;
      RECT 208.75 10.27 208.91 11.72 ;
      RECT 209.71 12 209.87 12.84 ;
      RECT 209.43 12 209.87 12.16 ;
      RECT 209.43 11.88 209.59 12.16 ;
      RECT 208.35 28.04 208.67 28.32 ;
      RECT 208.51 25.99 208.67 28.32 ;
      RECT 209.7 27.02 209.86 27.7 ;
      RECT 208.51 27.02 209.86 27.18 ;
      RECT 208.51 25.99 208.89 26.23 ;
      RECT 208.73 25.16 208.89 26.23 ;
      RECT 209.31 55.68 209.47 56.51 ;
      RECT 209.07 55.68 209.47 55.84 ;
      RECT 209.07 53.67 209.23 55.84 ;
      RECT 209.07 53.67 209.71 53.83 ;
      RECT 209.43 53.35 209.71 53.83 ;
      RECT 209.17 51.7 209.55 51.92 ;
      RECT 209.39 50.98 209.55 51.92 ;
      RECT 208.75 52.58 209.51 52.86 ;
      RECT 209.35 52.18 209.51 52.86 ;
      RECT 208.75 51.64 208.91 52.86 ;
      RECT 207.57 8.5 207.73 11.72 ;
      RECT 206.61 8.12 206.77 11.72 ;
      RECT 205.65 9.28 205.81 11.72 ;
      RECT 209.23 9.63 209.39 11.4 ;
      RECT 207.57 9.95 209.39 10.11 ;
      RECT 208.54 9.79 208.7 10.11 ;
      RECT 205.57 8.12 205.77 9.84 ;
      RECT 208.94 9.63 209.45 9.79 ;
      RECT 205.57 9.28 206.77 9.44 ;
      RECT 207.46 8.5 207.77 8.78 ;
      RECT 206.61 8.56 207.77 8.72 ;
      RECT 209.07 62.9 209.23 67.89 ;
      RECT 209.07 65.82 209.29 66.55 ;
      RECT 208.06 8.96 208.22 9.79 ;
      RECT 208.06 8.96 209.25 9.12 ;
      RECT 208.75 47.39 208.91 49.72 ;
      RECT 208.75 47.39 209.23 47.55 ;
      RECT 209.07 43.85 209.23 47.55 ;
      RECT 208.45 43.85 209.23 44.01 ;
      RECT 208.45 39.56 208.61 44.01 ;
      RECT 208.45 39.56 208.79 39.84 ;
      RECT 208.63 39.16 208.79 39.84 ;
      RECT 209.05 22.01 209.21 23.37 ;
      RECT 208.43 22.01 209.21 22.17 ;
      RECT 208.73 24.72 209.11 24.96 ;
      RECT 208.73 22.35 208.89 24.96 ;
      RECT 208.77 34.44 209.11 34.72 ;
      RECT 208.95 32.44 209.11 34.72 ;
      RECT 208.77 33.11 209.11 33.39 ;
      RECT 208.77 32.44 209.11 32.72 ;
      RECT 208.77 40.7 209.11 40.98 ;
      RECT 208.95 38.7 209.11 40.98 ;
      RECT 208.77 40.03 209.11 40.31 ;
      RECT 208.77 38.7 209.11 38.98 ;
      RECT 208.93 14.44 209.09 15.64 ;
      RECT 208.59 14.44 209.09 14.6 ;
      RECT 208.75 12.21 208.91 13.28 ;
      RECT 207.33 12.21 208.91 12.37 ;
      RECT 208.29 11.47 208.45 12.37 ;
      RECT 208.23 10.85 208.39 11.63 ;
      RECT 208.59 62.9 208.75 67.89 ;
      RECT 208.59 64.59 208.87 65.31 ;
      RECT 208.11 46.75 208.27 47.43 ;
      RECT 207.79 46.75 208.59 46.91 ;
      RECT 208.43 44.23 208.59 46.91 ;
      RECT 207.79 44.23 207.95 46.91 ;
      RECT 207.91 10.51 208.07 11.24 ;
      RECT 207.91 10.51 208.57 10.67 ;
      RECT 208.27 20.63 208.55 20.79 ;
      RECT 208.27 19.59 208.43 20.79 ;
      RECT 207.17 12.53 207.33 13.61 ;
      RECT 207.01 11.88 207.17 12.69 ;
      RECT 207.89 11.77 208.13 12.05 ;
      RECT 207.01 11.88 208.13 12.04 ;
      RECT 207.09 8.88 207.25 12.04 ;
      RECT 205.89 34.88 208.09 35.04 ;
      RECT 207.81 34.59 208.09 35.04 ;
      RECT 206.87 34.59 207.11 35.04 ;
      RECT 205.89 34.59 206.17 35.04 ;
      RECT 206.87 38.38 207.11 39.02 ;
      RECT 207.81 38.38 208.09 38.83 ;
      RECT 205.89 38.38 206.17 38.83 ;
      RECT 205.89 38.38 208.09 38.54 ;
      RECT 207.71 28.04 208.03 28.32 ;
      RECT 207.71 25.99 207.87 28.32 ;
      RECT 206.52 27.02 206.68 27.7 ;
      RECT 206.52 27.02 207.87 27.18 ;
      RECT 207.49 25.99 207.87 26.23 ;
      RECT 207.49 25.16 207.65 26.23 ;
      RECT 206.05 36.47 207.93 36.63 ;
      RECT 207.77 35.88 207.93 36.63 ;
      RECT 206.91 35.23 207.07 36.63 ;
      RECT 206.05 35.88 206.21 36.63 ;
      RECT 207.87 35.23 208.03 36.06 ;
      RECT 205.95 35.23 206.11 36.06 ;
      RECT 207.87 37.11 208.03 38.19 ;
      RECT 206.91 36.79 207.07 38.19 ;
      RECT 205.95 37.11 206.11 38.19 ;
      RECT 207.77 36.79 207.93 37.39 ;
      RECT 206.05 36.79 206.21 37.39 ;
      RECT 206.05 36.79 207.93 36.95 ;
      RECT 207.85 20.26 208.01 21.05 ;
      RECT 207.28 20.26 208.01 20.44 ;
      RECT 207.28 19.89 207.44 20.44 ;
      RECT 206.62 19.89 207.44 20.05 ;
      RECT 206.62 19.61 206.81 20.05 ;
      RECT 206.53 19.61 206.81 19.77 ;
      RECT 207.17 22.01 207.33 23.37 ;
      RECT 207.17 22.01 207.95 22.17 ;
      RECT 206.13 68.07 207.95 68.23 ;
      RECT 206.13 62.02 206.29 68.23 ;
      RECT 206.13 62.02 206.51 62.18 ;
      RECT 206.35 57.45 206.51 62.18 ;
      RECT 206.35 57.45 207.95 57.61 ;
      RECT 207.63 57.39 207.95 57.61 ;
      RECT 207.63 53.74 207.79 57.61 ;
      RECT 207.79 51.32 207.95 53.9 ;
      RECT 207.47 51.32 207.95 51.48 ;
      RECT 207.47 49.88 207.63 51.48 ;
      RECT 207.15 49.88 207.63 50.04 ;
      RECT 207.15 47.71 207.31 50.04 ;
      RECT 206.69 47.71 207.31 47.99 ;
      RECT 207.47 47.39 207.63 49.72 ;
      RECT 207.15 47.39 207.63 47.55 ;
      RECT 207.15 43.85 207.31 47.55 ;
      RECT 207.15 43.85 207.93 44.01 ;
      RECT 207.77 39.56 207.93 44.01 ;
      RECT 207.59 39.56 207.93 39.84 ;
      RECT 207.59 39.16 207.75 39.84 ;
      RECT 207.63 62.9 207.79 67.89 ;
      RECT 207.51 64.59 207.79 65.31 ;
      RECT 207.27 24.72 207.65 24.96 ;
      RECT 207.49 22.35 207.65 24.96 ;
      RECT 206.87 52.58 207.63 52.86 ;
      RECT 207.47 51.64 207.63 52.86 ;
      RECT 206.87 52.18 207.03 52.86 ;
      RECT 207.27 34.44 207.61 34.72 ;
      RECT 207.27 32.44 207.43 34.72 ;
      RECT 207.27 33.11 207.61 33.39 ;
      RECT 207.27 32.44 207.61 32.72 ;
      RECT 207.27 40.7 207.61 40.98 ;
      RECT 207.27 38.7 207.43 40.98 ;
      RECT 207.27 40.03 207.61 40.31 ;
      RECT 207.27 38.7 207.61 38.98 ;
      RECT 207.33 53.23 207.61 53.51 ;
      RECT 207.33 53.03 207.49 53.51 ;
      RECT 206.51 53.03 207.49 53.19 ;
      RECT 206.51 50.98 206.67 53.19 ;
      RECT 206.47 52.54 206.67 52.82 ;
      RECT 206.13 50.98 206.67 51.14 ;
      RECT 206.13 50.8 206.35 51.14 ;
      RECT 206.03 56.67 206.19 61.86 ;
      RECT 206.03 56.67 207.47 56.83 ;
      RECT 207.31 56 207.47 56.83 ;
      RECT 206.19 54.4 206.35 56.83 ;
      RECT 207.17 26.36 207.33 26.72 ;
      RECT 205.03 26.36 207.33 26.52 ;
      RECT 205.03 26.04 205.19 26.52 ;
      RECT 204.38 26.04 205.19 26.2 ;
      RECT 207.15 50.66 207.31 51.5 ;
      RECT 206.51 50.66 207.31 50.82 ;
      RECT 206.51 50.18 206.67 50.82 ;
      RECT 206.03 50.18 206.67 50.5 ;
      RECT 206.03 47.07 206.19 50.5 ;
      RECT 206.03 47.07 206.51 47.23 ;
      RECT 206.35 45.44 206.51 47.23 ;
      RECT 206.91 55.68 207.07 56.51 ;
      RECT 206.91 55.68 207.31 55.84 ;
      RECT 207.15 53.67 207.31 55.84 ;
      RECT 206.67 53.67 207.31 53.83 ;
      RECT 206.67 53.35 206.95 53.83 ;
      RECT 207.15 62.9 207.31 67.89 ;
      RECT 207.09 65.82 207.31 66.55 ;
      RECT 206.83 51.7 207.21 51.92 ;
      RECT 206.83 50.98 206.99 51.92 ;
      RECT 205 28.01 207.16 28.17 ;
      RECT 207 27.34 207.16 28.17 ;
      RECT 206.84 27.93 207.16 28.17 ;
      RECT 206 26.97 206.16 28.17 ;
      RECT 205 26.68 205.16 28.17 ;
      RECT 206.35 47.39 206.51 49.72 ;
      RECT 206.35 47.39 206.83 47.55 ;
      RECT 206.67 43.85 206.83 47.55 ;
      RECT 206.05 43.85 206.83 44.01 ;
      RECT 206.05 39.56 206.21 44.01 ;
      RECT 206.05 39.56 206.39 39.84 ;
      RECT 206.23 39.16 206.39 39.84 ;
      RECT 206.51 24.79 206.71 25.35 ;
      RECT 206.39 24.79 206.71 25.03 ;
      RECT 206.37 34.44 206.71 34.72 ;
      RECT 206.55 32.44 206.71 34.72 ;
      RECT 206.37 33.11 206.71 33.39 ;
      RECT 206.37 32.44 206.71 32.72 ;
      RECT 206.37 40.7 206.71 40.98 ;
      RECT 206.55 38.7 206.71 40.98 ;
      RECT 206.37 40.03 206.71 40.31 ;
      RECT 206.37 38.7 206.71 38.98 ;
      RECT 206.39 21.85 206.55 24.3 ;
      RECT 206.39 21.85 206.69 22.13 ;
      RECT 206.51 54.06 206.67 56.51 ;
      RECT 206.15 54.06 206.67 54.22 ;
      RECT 206.15 52.98 206.35 54.22 ;
      RECT 206.15 51.34 206.31 54.22 ;
      RECT 206.15 51.34 206.35 52.12 ;
      RECT 206.21 12.56 206.37 13.61 ;
      RECT 206.31 11.9 206.47 13.24 ;
      RECT 205.19 11.9 206.47 12.06 ;
      RECT 206.13 9.6 206.29 12.06 ;
      RECT 204.78 18.3 205.72 18.46 ;
      RECT 204.78 17.05 205.14 18.46 ;
      RECT 204.98 16.2 205.14 18.46 ;
      RECT 204.93 16.2 205.89 16.36 ;
      RECT 205.66 16.07 206.33 16.23 ;
      RECT 204.93 16.08 205.09 16.36 ;
      RECT 205.97 8.96 206.29 9.12 ;
      RECT 206.13 7.8 206.29 9.12 ;
      RECT 203.79 7.91 203.95 8.8 ;
      RECT 203.79 7.91 204.87 8.07 ;
      RECT 204.71 7.8 206.29 7.96 ;
      RECT 205.3 16.52 205.48 16.84 ;
      RECT 205.3 16.52 206.2 16.68 ;
      RECT 205.71 46.75 205.87 47.43 ;
      RECT 205.39 46.75 206.19 46.91 ;
      RECT 206.03 44.23 206.19 46.91 ;
      RECT 205.39 44.23 205.55 46.91 ;
      RECT 205.78 16.92 205.94 18.12 ;
      RECT 205.78 16.92 206.18 17.08 ;
      RECT 204.63 11.5 204.79 13.22 ;
      RECT 204.63 12.22 206.15 12.38 ;
      RECT 204.63 11.5 205.05 11.66 ;
      RECT 205.55 26.02 206.11 26.18 ;
      RECT 205.55 25.58 205.71 26.18 ;
      RECT 205.01 25.58 205.71 25.74 ;
      RECT 205.01 24 205.21 25.74 ;
      RECT 204.21 24.3 205.21 24.46 ;
      RECT 205.01 22.71 205.17 25.74 ;
      RECT 205.11 22.04 205.27 22.99 ;
      RECT 205.27 21.85 205.43 22.32 ;
      RECT 204.59 22.13 204.95 22.41 ;
      RECT 204.79 21.53 204.95 22.41 ;
      RECT 205.66 21.53 205.82 21.92 ;
      RECT 204.79 21.53 205.82 21.69 ;
      RECT 205.48 20.21 205.64 21.69 ;
      RECT 205.52 26.69 205.68 27.85 ;
      RECT 205.48 26.69 205.72 27.33 ;
      RECT 203.49 34.88 205.69 35.04 ;
      RECT 205.41 34.59 205.69 35.04 ;
      RECT 204.47 34.59 204.71 35.04 ;
      RECT 203.49 34.59 203.77 35.04 ;
      RECT 204.47 38.38 204.71 39.02 ;
      RECT 205.41 38.38 205.69 38.83 ;
      RECT 203.49 38.38 203.77 38.83 ;
      RECT 203.49 38.38 205.69 38.54 ;
      RECT 205.33 23.18 205.49 23.84 ;
      RECT 205.33 23.18 205.66 23.34 ;
      RECT 205.5 22.65 205.66 23.34 ;
      RECT 203.65 36.47 205.53 36.63 ;
      RECT 205.37 35.86 205.53 36.63 ;
      RECT 204.51 35.23 204.67 36.63 ;
      RECT 203.65 35.86 203.81 36.63 ;
      RECT 205.47 35.23 205.63 36.05 ;
      RECT 203.55 35.23 203.71 36.05 ;
      RECT 205.47 37.11 205.63 38.19 ;
      RECT 204.51 36.79 204.67 38.19 ;
      RECT 203.55 37.11 203.71 38.19 ;
      RECT 205.37 36.79 205.53 37.39 ;
      RECT 203.65 36.79 203.81 37.39 ;
      RECT 203.65 36.79 205.53 36.95 ;
      RECT 204.27 50.66 204.43 51.5 ;
      RECT 204.27 50.66 205.07 50.82 ;
      RECT 204.91 50.18 205.07 50.82 ;
      RECT 204.91 50.18 205.55 50.5 ;
      RECT 205.39 47.07 205.55 50.5 ;
      RECT 205.07 47.07 205.55 47.23 ;
      RECT 205.07 45.44 205.23 47.23 ;
      RECT 205.39 56.67 205.55 61.86 ;
      RECT 204.11 56.67 205.55 56.83 ;
      RECT 205.23 54.4 205.39 56.83 ;
      RECT 204.11 56 204.27 56.83 ;
      RECT 205.07 47.39 205.23 49.72 ;
      RECT 204.75 47.39 205.23 47.55 ;
      RECT 204.75 43.85 204.91 47.55 ;
      RECT 204.75 43.85 205.53 44.01 ;
      RECT 205.37 39.56 205.53 44.01 ;
      RECT 205.19 39.56 205.53 39.84 ;
      RECT 205.19 39.16 205.35 39.84 ;
      RECT 203.98 28.52 205.07 28.68 ;
      RECT 204.79 28.35 205.07 28.68 ;
      RECT 204.79 28.35 205.47 28.51 ;
      RECT 203.97 53.23 204.25 53.51 ;
      RECT 204.09 53.03 204.25 53.51 ;
      RECT 204.09 53.03 205.07 53.19 ;
      RECT 204.91 50.98 205.07 53.19 ;
      RECT 204.91 52.54 205.11 52.82 ;
      RECT 204.91 50.98 205.45 51.14 ;
      RECT 205.23 50.8 205.45 51.14 ;
      RECT 203.63 68.07 205.45 68.23 ;
      RECT 205.29 62.02 205.45 68.23 ;
      RECT 205.07 62.02 205.45 62.18 ;
      RECT 205.07 57.45 205.23 62.18 ;
      RECT 203.63 57.45 205.23 57.61 ;
      RECT 203.63 57.39 203.95 57.61 ;
      RECT 203.79 53.74 203.95 57.61 ;
      RECT 203.63 51.32 203.79 53.9 ;
      RECT 203.63 51.32 204.11 51.48 ;
      RECT 203.95 49.88 204.11 51.48 ;
      RECT 203.95 49.88 204.43 50.04 ;
      RECT 204.27 47.71 204.43 50.04 ;
      RECT 204.27 47.71 204.89 47.99 ;
      RECT 204.91 54.06 205.07 56.51 ;
      RECT 204.91 54.06 205.43 54.22 ;
      RECT 205.27 51.34 205.43 54.22 ;
      RECT 205.23 52.98 205.43 54.22 ;
      RECT 205.23 51.34 205.43 52.12 ;
      RECT 204.11 12.92 204.27 13.67 ;
      RECT 204.11 12.92 204.47 13.08 ;
      RECT 204.31 9.68 204.47 13.08 ;
      RECT 204.27 9.68 204.47 11.89 ;
      RECT 204.27 9.68 205.25 9.84 ;
      RECT 205.09 8.6 205.25 9.84 ;
      RECT 204.87 34.44 205.21 34.72 ;
      RECT 204.87 32.44 205.03 34.72 ;
      RECT 204.87 33.11 205.21 33.39 ;
      RECT 204.87 32.44 205.21 32.72 ;
      RECT 204.87 40.7 205.21 40.98 ;
      RECT 204.87 38.7 205.03 40.98 ;
      RECT 204.87 40.03 205.21 40.31 ;
      RECT 204.87 38.7 205.21 38.98 ;
      RECT 204.51 55.68 204.67 56.51 ;
      RECT 204.27 55.68 204.67 55.84 ;
      RECT 204.27 53.67 204.43 55.84 ;
      RECT 204.27 53.67 204.91 53.83 ;
      RECT 204.63 53.35 204.91 53.83 ;
      RECT 204.46 16.52 204.62 18.9 ;
      RECT 204.46 16.52 204.82 16.8 ;
      RECT 204.59 15.31 204.75 16.8 ;
      RECT 204.06 24.79 204.22 28.32 ;
      RECT 204.06 25.16 204.75 25.32 ;
      RECT 204.37 51.7 204.75 51.92 ;
      RECT 204.59 50.98 204.75 51.92 ;
      RECT 203.95 52.58 204.71 52.86 ;
      RECT 204.55 52.18 204.71 52.86 ;
      RECT 203.95 51.64 204.11 52.86 ;
      RECT 203.79 23.98 203.97 24.52 ;
      RECT 203.79 23.98 204.49 24.14 ;
      RECT 204.33 23.27 204.49 24.14 ;
      RECT 204.27 21.78 204.43 23.43 ;
      RECT 204.41 21.21 204.57 21.94 ;
      RECT 204.54 20.95 204.7 21.37 ;
      RECT 203.31 7.5 203.47 8.72 ;
      RECT 203.31 7.58 203.52 7.9 ;
      RECT 203.31 7.59 204.55 7.75 ;
      RECT 203.31 7.58 203.59 7.75 ;
      RECT 204.27 62.9 204.43 67.89 ;
      RECT 204.27 65.82 204.49 66.55 ;
      RECT 203.95 47.39 204.11 49.72 ;
      RECT 203.95 47.39 204.43 47.55 ;
      RECT 204.27 43.85 204.43 47.55 ;
      RECT 203.65 43.85 204.43 44.01 ;
      RECT 203.65 39.56 203.81 44.01 ;
      RECT 203.65 39.56 203.99 39.84 ;
      RECT 203.83 39.16 203.99 39.84 ;
      RECT 203.97 34.44 204.31 34.72 ;
      RECT 204.15 32.44 204.31 34.72 ;
      RECT 203.97 33.11 204.31 33.39 ;
      RECT 203.97 32.44 204.31 32.72 ;
      RECT 203.97 40.7 204.31 40.98 ;
      RECT 204.15 38.7 204.31 40.98 ;
      RECT 203.97 40.03 204.31 40.31 ;
      RECT 203.97 38.7 204.31 38.98 ;
      RECT 203.54 15.57 203.7 17.28 ;
      RECT 204.14 16.43 204.3 16.71 ;
      RECT 203.54 16.43 204.3 16.59 ;
      RECT 203.48 15.57 203.76 15.73 ;
      RECT 203.98 17.18 204.14 18.9 ;
      RECT 203.31 17.96 204.14 18.12 ;
      RECT 203.31 17.84 203.47 18.12 ;
      RECT 204.02 17.06 204.18 17.34 ;
      RECT 203.63 23.66 204.17 23.82 ;
      RECT 203.63 20.12 203.79 23.82 ;
      RECT 203.63 23.22 204.09 23.38 ;
      RECT 203.54 20.83 203.79 21.11 ;
      RECT 203.63 20.12 204.06 20.28 ;
      RECT 203.79 62.9 203.95 67.89 ;
      RECT 203.79 64.59 204.07 65.31 ;
      RECT 203.83 10.08 203.99 11.89 ;
      RECT 203.25 10.08 203.99 10.24 ;
      RECT 203.31 8.88 203.47 10.24 ;
      RECT 203.31 46.75 203.47 47.43 ;
      RECT 202.99 46.75 203.79 46.91 ;
      RECT 203.63 44.23 203.79 46.91 ;
      RECT 202.99 44.23 203.15 46.91 ;
      RECT 203.58 26.15 203.74 28.96 ;
      RECT 203.55 26.15 203.74 26.51 ;
      RECT 201.09 34.88 203.29 35.04 ;
      RECT 203.01 34.59 203.29 35.04 ;
      RECT 202.07 34.59 202.31 35.04 ;
      RECT 201.09 34.59 201.37 35.04 ;
      RECT 202.07 38.38 202.31 39.02 ;
      RECT 203.01 38.38 203.29 38.83 ;
      RECT 201.09 38.38 201.37 38.83 ;
      RECT 201.09 38.38 203.29 38.54 ;
      RECT 201.25 36.47 203.13 36.63 ;
      RECT 202.97 35.88 203.13 36.63 ;
      RECT 202.11 35.23 202.27 36.63 ;
      RECT 201.25 35.88 201.41 36.63 ;
      RECT 203.07 35.23 203.23 36.06 ;
      RECT 201.15 35.23 201.31 36.06 ;
      RECT 203.07 37.11 203.23 38.19 ;
      RECT 202.11 36.79 202.27 38.19 ;
      RECT 201.15 37.11 201.31 38.19 ;
      RECT 202.97 36.79 203.13 37.39 ;
      RECT 201.25 36.79 201.41 37.39 ;
      RECT 201.25 36.79 203.13 36.95 ;
      RECT 201.33 68.07 203.15 68.23 ;
      RECT 201.33 62.02 201.49 68.23 ;
      RECT 201.33 62.02 201.71 62.18 ;
      RECT 201.55 57.45 201.71 62.18 ;
      RECT 201.55 57.45 203.15 57.61 ;
      RECT 202.83 57.39 203.15 57.61 ;
      RECT 202.83 53.74 202.99 57.61 ;
      RECT 202.99 51.32 203.15 53.9 ;
      RECT 202.67 51.32 203.15 51.48 ;
      RECT 202.67 49.88 202.83 51.48 ;
      RECT 202.35 49.88 202.83 50.04 ;
      RECT 202.35 47.71 202.51 50.04 ;
      RECT 201.89 47.71 202.51 47.99 ;
      RECT 202.67 47.39 202.83 49.72 ;
      RECT 202.35 47.39 202.83 47.55 ;
      RECT 202.35 43.85 202.51 47.55 ;
      RECT 202.35 43.85 203.13 44.01 ;
      RECT 202.97 39.56 203.13 44.01 ;
      RECT 202.79 39.56 203.13 39.84 ;
      RECT 202.79 39.16 202.95 39.84 ;
      RECT 202.83 62.9 202.99 67.89 ;
      RECT 202.71 64.59 202.99 65.31 ;
      RECT 202.07 52.58 202.83 52.86 ;
      RECT 202.67 51.64 202.83 52.86 ;
      RECT 202.07 52.18 202.23 52.86 ;
      RECT 202.47 34.44 202.81 34.72 ;
      RECT 202.47 32.44 202.63 34.72 ;
      RECT 202.47 33.11 202.81 33.39 ;
      RECT 202.47 32.44 202.81 32.72 ;
      RECT 202.47 40.7 202.81 40.98 ;
      RECT 202.47 38.7 202.63 40.98 ;
      RECT 202.47 40.03 202.81 40.31 ;
      RECT 202.47 38.7 202.81 38.98 ;
      RECT 202.53 53.23 202.81 53.51 ;
      RECT 202.53 53.03 202.69 53.51 ;
      RECT 201.71 53.03 202.69 53.19 ;
      RECT 201.71 50.98 201.87 53.19 ;
      RECT 201.67 52.54 201.87 52.82 ;
      RECT 201.33 50.98 201.87 51.14 ;
      RECT 201.33 50.8 201.55 51.14 ;
      RECT 201.23 56.67 201.39 61.86 ;
      RECT 201.23 56.67 202.67 56.83 ;
      RECT 202.51 56 202.67 56.83 ;
      RECT 201.39 54.4 201.55 56.83 ;
      RECT 194.67 12.95 202.51 13.55 ;
      RECT 201.91 8.34 202.51 13.55 ;
      RECT 194.67 8.34 195.27 13.55 ;
      RECT 194.67 8.34 202.51 8.88 ;
      RECT 194.67 26.87 202.51 27.47 ;
      RECT 201.91 18.71 202.51 27.47 ;
      RECT 194.67 18.71 195.27 27.47 ;
      RECT 194.67 24.41 202.51 25.01 ;
      RECT 194.67 18.71 202.51 19.31 ;
      RECT 202.35 50.66 202.51 51.5 ;
      RECT 201.71 50.66 202.51 50.82 ;
      RECT 201.71 50.18 201.87 50.82 ;
      RECT 201.23 50.18 201.87 50.5 ;
      RECT 201.23 47.07 201.39 50.5 ;
      RECT 201.23 47.07 201.71 47.23 ;
      RECT 201.55 45.44 201.71 47.23 ;
      RECT 202.11 55.68 202.27 56.51 ;
      RECT 202.11 55.68 202.51 55.84 ;
      RECT 202.35 53.67 202.51 55.84 ;
      RECT 201.87 53.67 202.51 53.83 ;
      RECT 201.87 53.35 202.15 53.83 ;
      RECT 202.35 62.9 202.51 67.89 ;
      RECT 202.29 65.82 202.51 66.55 ;
      RECT 202.03 51.7 202.41 51.92 ;
      RECT 202.03 50.98 202.19 51.92 ;
      RECT 201.55 47.39 201.71 49.72 ;
      RECT 201.55 47.39 202.03 47.55 ;
      RECT 201.87 43.85 202.03 47.55 ;
      RECT 201.25 43.85 202.03 44.01 ;
      RECT 201.25 39.56 201.41 44.01 ;
      RECT 201.25 39.56 201.59 39.84 ;
      RECT 201.43 39.16 201.59 39.84 ;
      RECT 201.57 34.44 201.91 34.72 ;
      RECT 201.75 32.44 201.91 34.72 ;
      RECT 201.57 33.11 201.91 33.39 ;
      RECT 201.57 32.44 201.91 32.72 ;
      RECT 201.57 40.7 201.91 40.98 ;
      RECT 201.75 38.7 201.91 40.98 ;
      RECT 201.57 40.03 201.91 40.31 ;
      RECT 201.57 38.7 201.91 38.98 ;
      RECT 201.71 54.06 201.87 56.51 ;
      RECT 201.35 54.06 201.87 54.22 ;
      RECT 201.35 52.98 201.55 54.22 ;
      RECT 201.35 51.34 201.51 54.22 ;
      RECT 201.35 51.34 201.55 52.12 ;
      RECT 200.91 46.75 201.07 47.43 ;
      RECT 200.59 46.75 201.39 46.91 ;
      RECT 201.23 44.23 201.39 46.91 ;
      RECT 200.59 44.23 200.75 46.91 ;
      RECT 198.69 34.88 200.89 35.04 ;
      RECT 200.61 34.59 200.89 35.04 ;
      RECT 199.67 34.59 199.91 35.04 ;
      RECT 198.69 34.59 198.97 35.04 ;
      RECT 199.67 38.38 199.91 39.02 ;
      RECT 200.61 38.38 200.89 38.83 ;
      RECT 198.69 38.38 198.97 38.83 ;
      RECT 198.69 38.38 200.89 38.54 ;
      RECT 198.85 36.47 200.73 36.63 ;
      RECT 200.57 35.86 200.73 36.63 ;
      RECT 199.71 35.23 199.87 36.63 ;
      RECT 198.85 35.86 199.01 36.63 ;
      RECT 200.67 35.23 200.83 36.05 ;
      RECT 198.75 35.23 198.91 36.05 ;
      RECT 200.67 37.11 200.83 38.19 ;
      RECT 199.71 36.79 199.87 38.19 ;
      RECT 198.75 37.11 198.91 38.19 ;
      RECT 200.57 36.79 200.73 37.39 ;
      RECT 198.85 36.79 199.01 37.39 ;
      RECT 198.85 36.79 200.73 36.95 ;
      RECT 199.47 50.66 199.63 51.5 ;
      RECT 199.47 50.66 200.27 50.82 ;
      RECT 200.11 50.18 200.27 50.82 ;
      RECT 200.11 50.18 200.75 50.5 ;
      RECT 200.59 47.07 200.75 50.5 ;
      RECT 200.27 47.07 200.75 47.23 ;
      RECT 200.27 45.44 200.43 47.23 ;
      RECT 200.59 56.67 200.75 61.86 ;
      RECT 199.31 56.67 200.75 56.83 ;
      RECT 200.43 54.4 200.59 56.83 ;
      RECT 199.31 56 199.47 56.83 ;
      RECT 200.27 47.39 200.43 49.72 ;
      RECT 199.95 47.39 200.43 47.55 ;
      RECT 199.95 43.85 200.11 47.55 ;
      RECT 199.95 43.85 200.73 44.01 ;
      RECT 200.57 39.56 200.73 44.01 ;
      RECT 200.39 39.56 200.73 39.84 ;
      RECT 200.39 39.16 200.55 39.84 ;
      RECT 199.17 53.23 199.45 53.51 ;
      RECT 199.29 53.03 199.45 53.51 ;
      RECT 199.29 53.03 200.27 53.19 ;
      RECT 200.11 50.98 200.27 53.19 ;
      RECT 200.11 52.54 200.31 52.82 ;
      RECT 200.11 50.98 200.65 51.14 ;
      RECT 200.43 50.8 200.65 51.14 ;
      RECT 198.83 68.07 200.65 68.23 ;
      RECT 200.49 62.02 200.65 68.23 ;
      RECT 200.27 62.02 200.65 62.18 ;
      RECT 200.27 57.45 200.43 62.18 ;
      RECT 198.83 57.45 200.43 57.61 ;
      RECT 198.83 57.39 199.15 57.61 ;
      RECT 198.99 53.74 199.15 57.61 ;
      RECT 198.83 51.32 198.99 53.9 ;
      RECT 198.83 51.32 199.31 51.48 ;
      RECT 199.15 49.88 199.31 51.48 ;
      RECT 199.15 49.88 199.63 50.04 ;
      RECT 199.47 47.71 199.63 50.04 ;
      RECT 199.47 47.71 200.09 47.99 ;
      RECT 200.11 54.06 200.27 56.51 ;
      RECT 200.11 54.06 200.63 54.22 ;
      RECT 200.47 51.34 200.63 54.22 ;
      RECT 200.43 52.98 200.63 54.22 ;
      RECT 200.43 51.34 200.63 52.12 ;
      RECT 200.07 34.44 200.41 34.72 ;
      RECT 200.07 32.44 200.23 34.72 ;
      RECT 200.07 33.11 200.41 33.39 ;
      RECT 200.07 32.44 200.41 32.72 ;
      RECT 200.07 40.7 200.41 40.98 ;
      RECT 200.07 38.7 200.23 40.98 ;
      RECT 200.07 40.03 200.41 40.31 ;
      RECT 200.07 38.7 200.41 38.98 ;
      RECT 199.71 55.68 199.87 56.51 ;
      RECT 199.47 55.68 199.87 55.84 ;
      RECT 199.47 53.67 199.63 55.84 ;
      RECT 199.47 53.67 200.11 53.83 ;
      RECT 199.83 53.35 200.11 53.83 ;
      RECT 199.57 51.7 199.95 51.92 ;
      RECT 199.79 50.98 199.95 51.92 ;
      RECT 199.15 52.58 199.91 52.86 ;
      RECT 199.75 52.18 199.91 52.86 ;
      RECT 199.15 51.64 199.31 52.86 ;
      RECT 199.47 62.9 199.63 67.89 ;
      RECT 199.47 65.82 199.69 66.55 ;
      RECT 199.15 47.39 199.31 49.72 ;
      RECT 199.15 47.39 199.63 47.55 ;
      RECT 199.47 43.85 199.63 47.55 ;
      RECT 198.85 43.85 199.63 44.01 ;
      RECT 198.85 39.56 199.01 44.01 ;
      RECT 198.85 39.56 199.19 39.84 ;
      RECT 199.03 39.16 199.19 39.84 ;
      RECT 199.17 34.44 199.51 34.72 ;
      RECT 199.35 32.44 199.51 34.72 ;
      RECT 199.17 33.11 199.51 33.39 ;
      RECT 199.17 32.44 199.51 32.72 ;
      RECT 199.17 40.7 199.51 40.98 ;
      RECT 199.35 38.7 199.51 40.98 ;
      RECT 199.17 40.03 199.51 40.31 ;
      RECT 199.17 38.7 199.51 38.98 ;
      RECT 198.99 62.9 199.15 67.89 ;
      RECT 198.99 64.59 199.27 65.31 ;
      RECT 198.51 46.75 198.67 47.43 ;
      RECT 198.19 46.75 198.99 46.91 ;
      RECT 198.83 44.23 198.99 46.91 ;
      RECT 198.19 44.23 198.35 46.91 ;
      RECT 196.29 34.88 198.49 35.04 ;
      RECT 198.21 34.59 198.49 35.04 ;
      RECT 197.27 34.59 197.51 35.04 ;
      RECT 196.29 34.59 196.57 35.04 ;
      RECT 197.27 38.38 197.51 39.02 ;
      RECT 198.21 38.38 198.49 38.83 ;
      RECT 196.29 38.38 196.57 38.83 ;
      RECT 196.29 38.38 198.49 38.54 ;
      RECT 196.45 36.47 198.33 36.63 ;
      RECT 198.17 35.88 198.33 36.63 ;
      RECT 197.31 35.23 197.47 36.63 ;
      RECT 196.45 35.88 196.61 36.63 ;
      RECT 198.27 35.23 198.43 36.06 ;
      RECT 196.35 35.23 196.51 36.06 ;
      RECT 198.27 37.11 198.43 38.19 ;
      RECT 197.31 36.79 197.47 38.19 ;
      RECT 196.35 37.11 196.51 38.19 ;
      RECT 198.17 36.79 198.33 37.39 ;
      RECT 196.45 36.79 196.61 37.39 ;
      RECT 196.45 36.79 198.33 36.95 ;
      RECT 196.53 68.07 198.35 68.23 ;
      RECT 196.53 62.02 196.69 68.23 ;
      RECT 196.53 62.02 196.91 62.18 ;
      RECT 196.75 57.45 196.91 62.18 ;
      RECT 196.75 57.45 198.35 57.61 ;
      RECT 198.03 57.39 198.35 57.61 ;
      RECT 198.03 53.74 198.19 57.61 ;
      RECT 198.19 51.32 198.35 53.9 ;
      RECT 197.87 51.32 198.35 51.48 ;
      RECT 197.87 49.88 198.03 51.48 ;
      RECT 197.55 49.88 198.03 50.04 ;
      RECT 197.55 47.71 197.71 50.04 ;
      RECT 197.09 47.71 197.71 47.99 ;
      RECT 197.87 47.39 198.03 49.72 ;
      RECT 197.55 47.39 198.03 47.55 ;
      RECT 197.55 43.85 197.71 47.55 ;
      RECT 197.55 43.85 198.33 44.01 ;
      RECT 198.17 39.56 198.33 44.01 ;
      RECT 197.99 39.56 198.33 39.84 ;
      RECT 197.99 39.16 198.15 39.84 ;
      RECT 198.03 62.9 198.19 67.89 ;
      RECT 197.91 64.59 198.19 65.31 ;
      RECT 197.27 52.58 198.03 52.86 ;
      RECT 197.87 51.64 198.03 52.86 ;
      RECT 197.27 52.18 197.43 52.86 ;
      RECT 197.67 34.44 198.01 34.72 ;
      RECT 197.67 32.44 197.83 34.72 ;
      RECT 197.67 33.11 198.01 33.39 ;
      RECT 197.67 32.44 198.01 32.72 ;
      RECT 197.67 40.7 198.01 40.98 ;
      RECT 197.67 38.7 197.83 40.98 ;
      RECT 197.67 40.03 198.01 40.31 ;
      RECT 197.67 38.7 198.01 38.98 ;
      RECT 197.73 53.23 198.01 53.51 ;
      RECT 197.73 53.03 197.89 53.51 ;
      RECT 196.91 53.03 197.89 53.19 ;
      RECT 196.91 50.98 197.07 53.19 ;
      RECT 196.87 52.54 197.07 52.82 ;
      RECT 196.53 50.98 197.07 51.14 ;
      RECT 196.53 50.8 196.75 51.14 ;
      RECT 196.43 56.67 196.59 61.86 ;
      RECT 196.43 56.67 197.87 56.83 ;
      RECT 197.71 56 197.87 56.83 ;
      RECT 196.59 54.4 196.75 56.83 ;
      RECT 197.55 50.66 197.71 51.5 ;
      RECT 196.91 50.66 197.71 50.82 ;
      RECT 196.91 50.18 197.07 50.82 ;
      RECT 196.43 50.18 197.07 50.5 ;
      RECT 196.43 47.07 196.59 50.5 ;
      RECT 196.43 47.07 196.91 47.23 ;
      RECT 196.75 45.44 196.91 47.23 ;
      RECT 197.31 55.68 197.47 56.51 ;
      RECT 197.31 55.68 197.71 55.84 ;
      RECT 197.55 53.67 197.71 55.84 ;
      RECT 197.07 53.67 197.71 53.83 ;
      RECT 197.07 53.35 197.35 53.83 ;
      RECT 197.55 62.9 197.71 67.89 ;
      RECT 197.49 65.82 197.71 66.55 ;
      RECT 197.23 51.7 197.61 51.92 ;
      RECT 197.23 50.98 197.39 51.92 ;
      RECT 196.75 47.39 196.91 49.72 ;
      RECT 196.75 47.39 197.23 47.55 ;
      RECT 197.07 43.85 197.23 47.55 ;
      RECT 196.45 43.85 197.23 44.01 ;
      RECT 196.45 39.56 196.61 44.01 ;
      RECT 196.45 39.56 196.79 39.84 ;
      RECT 196.63 39.16 196.79 39.84 ;
      RECT 196.77 34.44 197.11 34.72 ;
      RECT 196.95 32.44 197.11 34.72 ;
      RECT 196.77 33.11 197.11 33.39 ;
      RECT 196.77 32.44 197.11 32.72 ;
      RECT 196.77 40.7 197.11 40.98 ;
      RECT 196.95 38.7 197.11 40.98 ;
      RECT 196.77 40.03 197.11 40.31 ;
      RECT 196.77 38.7 197.11 38.98 ;
      RECT 196.91 54.06 197.07 56.51 ;
      RECT 196.55 54.06 197.07 54.22 ;
      RECT 196.55 52.98 196.75 54.22 ;
      RECT 196.55 51.34 196.71 54.22 ;
      RECT 196.55 51.34 196.75 52.12 ;
      RECT 196.11 46.75 196.27 47.43 ;
      RECT 195.79 46.75 196.59 46.91 ;
      RECT 196.43 44.23 196.59 46.91 ;
      RECT 195.79 44.23 195.95 46.91 ;
      RECT 193.89 34.88 196.09 35.04 ;
      RECT 195.81 34.59 196.09 35.04 ;
      RECT 194.87 34.59 195.11 35.04 ;
      RECT 193.89 34.59 194.17 35.04 ;
      RECT 194.87 38.38 195.11 39.02 ;
      RECT 195.81 38.38 196.09 38.83 ;
      RECT 193.89 38.38 194.17 38.83 ;
      RECT 193.89 38.38 196.09 38.54 ;
      RECT 194.05 36.47 195.93 36.63 ;
      RECT 195.77 35.86 195.93 36.63 ;
      RECT 194.91 35.23 195.07 36.63 ;
      RECT 194.05 35.86 194.21 36.63 ;
      RECT 195.87 35.23 196.03 36.05 ;
      RECT 193.95 35.23 194.11 36.05 ;
      RECT 195.87 37.11 196.03 38.19 ;
      RECT 194.91 36.79 195.07 38.19 ;
      RECT 193.95 37.11 194.11 38.19 ;
      RECT 195.77 36.79 195.93 37.39 ;
      RECT 194.05 36.79 194.21 37.39 ;
      RECT 194.05 36.79 195.93 36.95 ;
      RECT 194.67 50.66 194.83 51.5 ;
      RECT 194.67 50.66 195.47 50.82 ;
      RECT 195.31 50.18 195.47 50.82 ;
      RECT 195.31 50.18 195.95 50.5 ;
      RECT 195.79 47.07 195.95 50.5 ;
      RECT 195.47 47.07 195.95 47.23 ;
      RECT 195.47 45.44 195.63 47.23 ;
      RECT 195.79 56.67 195.95 61.86 ;
      RECT 194.51 56.67 195.95 56.83 ;
      RECT 195.63 54.4 195.79 56.83 ;
      RECT 194.51 56 194.67 56.83 ;
      RECT 195.47 47.39 195.63 49.72 ;
      RECT 195.15 47.39 195.63 47.55 ;
      RECT 195.15 43.85 195.31 47.55 ;
      RECT 195.15 43.85 195.93 44.01 ;
      RECT 195.77 39.56 195.93 44.01 ;
      RECT 195.59 39.56 195.93 39.84 ;
      RECT 195.59 39.16 195.75 39.84 ;
      RECT 194.37 53.23 194.65 53.51 ;
      RECT 194.49 53.03 194.65 53.51 ;
      RECT 194.49 53.03 195.47 53.19 ;
      RECT 195.31 50.98 195.47 53.19 ;
      RECT 195.31 52.54 195.51 52.82 ;
      RECT 195.31 50.98 195.85 51.14 ;
      RECT 195.63 50.8 195.85 51.14 ;
      RECT 194.03 68.07 195.85 68.23 ;
      RECT 195.69 62.02 195.85 68.23 ;
      RECT 195.47 62.02 195.85 62.18 ;
      RECT 195.47 57.45 195.63 62.18 ;
      RECT 194.03 57.45 195.63 57.61 ;
      RECT 194.03 57.39 194.35 57.61 ;
      RECT 194.19 53.74 194.35 57.61 ;
      RECT 194.03 51.32 194.19 53.9 ;
      RECT 194.03 51.32 194.51 51.48 ;
      RECT 194.35 49.88 194.51 51.48 ;
      RECT 194.35 49.88 194.83 50.04 ;
      RECT 194.67 47.71 194.83 50.04 ;
      RECT 194.67 47.71 195.29 47.99 ;
      RECT 195.31 54.06 195.47 56.51 ;
      RECT 195.31 54.06 195.83 54.22 ;
      RECT 195.67 51.34 195.83 54.22 ;
      RECT 195.63 52.98 195.83 54.22 ;
      RECT 195.63 51.34 195.83 52.12 ;
      RECT 195.27 34.44 195.61 34.72 ;
      RECT 195.27 32.44 195.43 34.72 ;
      RECT 195.27 33.11 195.61 33.39 ;
      RECT 195.27 32.44 195.61 32.72 ;
      RECT 195.27 40.7 195.61 40.98 ;
      RECT 195.27 38.7 195.43 40.98 ;
      RECT 195.27 40.03 195.61 40.31 ;
      RECT 195.27 38.7 195.61 38.98 ;
      RECT 194.91 55.68 195.07 56.51 ;
      RECT 194.67 55.68 195.07 55.84 ;
      RECT 194.67 53.67 194.83 55.84 ;
      RECT 194.67 53.67 195.31 53.83 ;
      RECT 195.03 53.35 195.31 53.83 ;
      RECT 194.77 51.7 195.15 51.92 ;
      RECT 194.99 50.98 195.15 51.92 ;
      RECT 194.35 52.58 195.11 52.86 ;
      RECT 194.95 52.18 195.11 52.86 ;
      RECT 194.35 51.64 194.51 52.86 ;
      RECT 194.67 62.9 194.83 67.89 ;
      RECT 194.67 65.82 194.89 66.55 ;
      RECT 194.35 47.39 194.51 49.72 ;
      RECT 194.35 47.39 194.83 47.55 ;
      RECT 194.67 43.85 194.83 47.55 ;
      RECT 194.05 43.85 194.83 44.01 ;
      RECT 194.05 39.56 194.21 44.01 ;
      RECT 194.05 39.56 194.39 39.84 ;
      RECT 194.23 39.16 194.39 39.84 ;
      RECT 192.39 6.84 193.99 7.24 ;
      RECT 193.39 6.24 194.79 6.84 ;
      RECT 191.59 6.24 192.99 6.84 ;
      RECT 194.37 34.44 194.71 34.72 ;
      RECT 194.55 32.44 194.71 34.72 ;
      RECT 194.37 33.11 194.71 33.39 ;
      RECT 194.37 32.44 194.71 32.72 ;
      RECT 194.37 40.7 194.71 40.98 ;
      RECT 194.55 38.7 194.71 40.98 ;
      RECT 194.37 40.03 194.71 40.31 ;
      RECT 194.37 38.7 194.71 38.98 ;
      RECT 194.19 62.9 194.35 67.89 ;
      RECT 194.19 64.59 194.47 65.31 ;
      RECT 193.71 46.75 193.87 47.43 ;
      RECT 193.71 46.75 194.19 46.91 ;
      RECT 194.03 44.23 194.19 46.91 ;
      RECT 192.51 46.75 192.67 47.43 ;
      RECT 192.19 46.75 192.67 46.91 ;
      RECT 192.19 44.23 192.35 46.91 ;
      RECT 190.29 34.88 192.49 35.04 ;
      RECT 192.21 34.59 192.49 35.04 ;
      RECT 191.27 34.59 191.51 35.04 ;
      RECT 190.29 34.59 190.57 35.04 ;
      RECT 191.27 38.38 191.51 39.02 ;
      RECT 192.21 38.38 192.49 38.83 ;
      RECT 190.29 38.38 190.57 38.83 ;
      RECT 190.29 38.38 192.49 38.54 ;
      RECT 190.45 36.47 192.33 36.63 ;
      RECT 192.17 35.88 192.33 36.63 ;
      RECT 191.31 35.23 191.47 36.63 ;
      RECT 190.45 35.88 190.61 36.63 ;
      RECT 192.27 35.23 192.43 36.06 ;
      RECT 190.35 35.23 190.51 36.06 ;
      RECT 192.27 37.11 192.43 38.19 ;
      RECT 191.31 36.79 191.47 38.19 ;
      RECT 190.35 37.11 190.51 38.19 ;
      RECT 192.17 36.79 192.33 37.39 ;
      RECT 190.45 36.79 190.61 37.39 ;
      RECT 190.45 36.79 192.33 36.95 ;
      RECT 190.53 68.07 192.35 68.23 ;
      RECT 190.53 62.02 190.69 68.23 ;
      RECT 190.53 62.02 190.91 62.18 ;
      RECT 190.75 57.45 190.91 62.18 ;
      RECT 190.75 57.45 192.35 57.61 ;
      RECT 192.03 57.39 192.35 57.61 ;
      RECT 192.03 53.74 192.19 57.61 ;
      RECT 192.19 51.32 192.35 53.9 ;
      RECT 191.87 51.32 192.35 51.48 ;
      RECT 191.87 49.88 192.03 51.48 ;
      RECT 191.55 49.88 192.03 50.04 ;
      RECT 191.55 47.71 191.71 50.04 ;
      RECT 191.09 47.71 191.71 47.99 ;
      RECT 191.87 47.39 192.03 49.72 ;
      RECT 191.55 47.39 192.03 47.55 ;
      RECT 191.55 43.85 191.71 47.55 ;
      RECT 191.55 43.85 192.33 44.01 ;
      RECT 192.17 39.56 192.33 44.01 ;
      RECT 191.99 39.56 192.33 39.84 ;
      RECT 191.99 39.16 192.15 39.84 ;
      RECT 192.03 62.9 192.19 67.89 ;
      RECT 191.91 64.59 192.19 65.31 ;
      RECT 191.27 52.58 192.03 52.86 ;
      RECT 191.87 51.64 192.03 52.86 ;
      RECT 191.27 52.18 191.43 52.86 ;
      RECT 191.67 34.44 192.01 34.72 ;
      RECT 191.67 32.44 191.83 34.72 ;
      RECT 191.67 33.11 192.01 33.39 ;
      RECT 191.67 32.44 192.01 32.72 ;
      RECT 191.67 40.7 192.01 40.98 ;
      RECT 191.67 38.7 191.83 40.98 ;
      RECT 191.67 40.03 192.01 40.31 ;
      RECT 191.67 38.7 192.01 38.98 ;
      RECT 191.73 53.23 192.01 53.51 ;
      RECT 191.73 53.03 191.89 53.51 ;
      RECT 190.91 53.03 191.89 53.19 ;
      RECT 190.91 50.98 191.07 53.19 ;
      RECT 190.87 52.54 191.07 52.82 ;
      RECT 190.53 50.98 191.07 51.14 ;
      RECT 190.53 50.8 190.75 51.14 ;
      RECT 190.43 56.67 190.59 61.86 ;
      RECT 190.43 56.67 191.87 56.83 ;
      RECT 191.71 56 191.87 56.83 ;
      RECT 190.59 54.4 190.75 56.83 ;
      RECT 183.87 12.95 191.71 13.55 ;
      RECT 191.11 8.34 191.71 13.55 ;
      RECT 183.87 8.34 184.47 13.55 ;
      RECT 183.87 8.34 191.71 8.88 ;
      RECT 183.87 26.87 191.71 27.47 ;
      RECT 191.11 18.71 191.71 27.47 ;
      RECT 183.87 18.71 184.47 27.47 ;
      RECT 183.87 24.41 191.71 25.01 ;
      RECT 183.87 18.71 191.71 19.31 ;
      RECT 191.55 50.66 191.71 51.5 ;
      RECT 190.91 50.66 191.71 50.82 ;
      RECT 190.91 50.18 191.07 50.82 ;
      RECT 190.43 50.18 191.07 50.5 ;
      RECT 190.43 47.07 190.59 50.5 ;
      RECT 190.43 47.07 190.91 47.23 ;
      RECT 190.75 45.44 190.91 47.23 ;
      RECT 191.31 55.68 191.47 56.51 ;
      RECT 191.31 55.68 191.71 55.84 ;
      RECT 191.55 53.67 191.71 55.84 ;
      RECT 191.07 53.67 191.71 53.83 ;
      RECT 191.07 53.35 191.35 53.83 ;
      RECT 191.55 62.9 191.71 67.89 ;
      RECT 191.49 65.82 191.71 66.55 ;
      RECT 191.23 51.7 191.61 51.92 ;
      RECT 191.23 50.98 191.39 51.92 ;
      RECT 190.75 47.39 190.91 49.72 ;
      RECT 190.75 47.39 191.23 47.55 ;
      RECT 191.07 43.85 191.23 47.55 ;
      RECT 190.45 43.85 191.23 44.01 ;
      RECT 190.45 39.56 190.61 44.01 ;
      RECT 190.45 39.56 190.79 39.84 ;
      RECT 190.63 39.16 190.79 39.84 ;
      RECT 190.77 34.44 191.11 34.72 ;
      RECT 190.95 32.44 191.11 34.72 ;
      RECT 190.77 33.11 191.11 33.39 ;
      RECT 190.77 32.44 191.11 32.72 ;
      RECT 190.77 40.7 191.11 40.98 ;
      RECT 190.95 38.7 191.11 40.98 ;
      RECT 190.77 40.03 191.11 40.31 ;
      RECT 190.77 38.7 191.11 38.98 ;
      RECT 190.91 54.06 191.07 56.51 ;
      RECT 190.55 54.06 191.07 54.22 ;
      RECT 190.55 52.98 190.75 54.22 ;
      RECT 190.55 51.34 190.71 54.22 ;
      RECT 190.55 51.34 190.75 52.12 ;
      RECT 190.11 46.75 190.27 47.43 ;
      RECT 189.79 46.75 190.59 46.91 ;
      RECT 190.43 44.23 190.59 46.91 ;
      RECT 189.79 44.23 189.95 46.91 ;
      RECT 187.89 34.88 190.09 35.04 ;
      RECT 189.81 34.59 190.09 35.04 ;
      RECT 188.87 34.59 189.11 35.04 ;
      RECT 187.89 34.59 188.17 35.04 ;
      RECT 188.87 38.38 189.11 39.02 ;
      RECT 189.81 38.38 190.09 38.83 ;
      RECT 187.89 38.38 188.17 38.83 ;
      RECT 187.89 38.38 190.09 38.54 ;
      RECT 188.05 36.47 189.93 36.63 ;
      RECT 189.77 35.86 189.93 36.63 ;
      RECT 188.91 35.23 189.07 36.63 ;
      RECT 188.05 35.86 188.21 36.63 ;
      RECT 189.87 35.23 190.03 36.05 ;
      RECT 187.95 35.23 188.11 36.05 ;
      RECT 189.87 37.11 190.03 38.19 ;
      RECT 188.91 36.79 189.07 38.19 ;
      RECT 187.95 37.11 188.11 38.19 ;
      RECT 189.77 36.79 189.93 37.39 ;
      RECT 188.05 36.79 188.21 37.39 ;
      RECT 188.05 36.79 189.93 36.95 ;
      RECT 188.67 50.66 188.83 51.5 ;
      RECT 188.67 50.66 189.47 50.82 ;
      RECT 189.31 50.18 189.47 50.82 ;
      RECT 189.31 50.18 189.95 50.5 ;
      RECT 189.79 47.07 189.95 50.5 ;
      RECT 189.47 47.07 189.95 47.23 ;
      RECT 189.47 45.44 189.63 47.23 ;
      RECT 189.79 56.67 189.95 61.86 ;
      RECT 188.51 56.67 189.95 56.83 ;
      RECT 189.63 54.4 189.79 56.83 ;
      RECT 188.51 56 188.67 56.83 ;
      RECT 189.47 47.39 189.63 49.72 ;
      RECT 189.15 47.39 189.63 47.55 ;
      RECT 189.15 43.85 189.31 47.55 ;
      RECT 189.15 43.85 189.93 44.01 ;
      RECT 189.77 39.56 189.93 44.01 ;
      RECT 189.59 39.56 189.93 39.84 ;
      RECT 189.59 39.16 189.75 39.84 ;
      RECT 188.37 53.23 188.65 53.51 ;
      RECT 188.49 53.03 188.65 53.51 ;
      RECT 188.49 53.03 189.47 53.19 ;
      RECT 189.31 50.98 189.47 53.19 ;
      RECT 189.31 52.54 189.51 52.82 ;
      RECT 189.31 50.98 189.85 51.14 ;
      RECT 189.63 50.8 189.85 51.14 ;
      RECT 188.03 68.07 189.85 68.23 ;
      RECT 189.69 62.02 189.85 68.23 ;
      RECT 189.47 62.02 189.85 62.18 ;
      RECT 189.47 57.45 189.63 62.18 ;
      RECT 188.03 57.45 189.63 57.61 ;
      RECT 188.03 57.39 188.35 57.61 ;
      RECT 188.19 53.74 188.35 57.61 ;
      RECT 188.03 51.32 188.19 53.9 ;
      RECT 188.03 51.32 188.51 51.48 ;
      RECT 188.35 49.88 188.51 51.48 ;
      RECT 188.35 49.88 188.83 50.04 ;
      RECT 188.67 47.71 188.83 50.04 ;
      RECT 188.67 47.71 189.29 47.99 ;
      RECT 189.31 54.06 189.47 56.51 ;
      RECT 189.31 54.06 189.83 54.22 ;
      RECT 189.67 51.34 189.83 54.22 ;
      RECT 189.63 52.98 189.83 54.22 ;
      RECT 189.63 51.34 189.83 52.12 ;
      RECT 189.27 34.44 189.61 34.72 ;
      RECT 189.27 32.44 189.43 34.72 ;
      RECT 189.27 33.11 189.61 33.39 ;
      RECT 189.27 32.44 189.61 32.72 ;
      RECT 189.27 40.7 189.61 40.98 ;
      RECT 189.27 38.7 189.43 40.98 ;
      RECT 189.27 40.03 189.61 40.31 ;
      RECT 189.27 38.7 189.61 38.98 ;
      RECT 188.91 55.68 189.07 56.51 ;
      RECT 188.67 55.68 189.07 55.84 ;
      RECT 188.67 53.67 188.83 55.84 ;
      RECT 188.67 53.67 189.31 53.83 ;
      RECT 189.03 53.35 189.31 53.83 ;
      RECT 188.77 51.7 189.15 51.92 ;
      RECT 188.99 50.98 189.15 51.92 ;
      RECT 188.35 52.58 189.11 52.86 ;
      RECT 188.95 52.18 189.11 52.86 ;
      RECT 188.35 51.64 188.51 52.86 ;
      RECT 188.67 62.9 188.83 67.89 ;
      RECT 188.67 65.82 188.89 66.55 ;
      RECT 188.35 47.39 188.51 49.72 ;
      RECT 188.35 47.39 188.83 47.55 ;
      RECT 188.67 43.85 188.83 47.55 ;
      RECT 188.05 43.85 188.83 44.01 ;
      RECT 188.05 39.56 188.21 44.01 ;
      RECT 188.05 39.56 188.39 39.84 ;
      RECT 188.23 39.16 188.39 39.84 ;
      RECT 188.37 34.44 188.71 34.72 ;
      RECT 188.55 32.44 188.71 34.72 ;
      RECT 188.37 33.11 188.71 33.39 ;
      RECT 188.37 32.44 188.71 32.72 ;
      RECT 188.37 40.7 188.71 40.98 ;
      RECT 188.55 38.7 188.71 40.98 ;
      RECT 188.37 40.03 188.71 40.31 ;
      RECT 188.37 38.7 188.71 38.98 ;
      RECT 188.19 62.9 188.35 67.89 ;
      RECT 188.19 64.59 188.47 65.31 ;
      RECT 187.71 46.75 187.87 47.43 ;
      RECT 187.39 46.75 188.19 46.91 ;
      RECT 188.03 44.23 188.19 46.91 ;
      RECT 187.39 44.23 187.55 46.91 ;
      RECT 185.49 34.88 187.69 35.04 ;
      RECT 187.41 34.59 187.69 35.04 ;
      RECT 186.47 34.59 186.71 35.04 ;
      RECT 185.49 34.59 185.77 35.04 ;
      RECT 186.47 38.38 186.71 39.02 ;
      RECT 187.41 38.38 187.69 38.83 ;
      RECT 185.49 38.38 185.77 38.83 ;
      RECT 185.49 38.38 187.69 38.54 ;
      RECT 185.65 36.47 187.53 36.63 ;
      RECT 187.37 35.88 187.53 36.63 ;
      RECT 186.51 35.23 186.67 36.63 ;
      RECT 185.65 35.88 185.81 36.63 ;
      RECT 187.47 35.23 187.63 36.06 ;
      RECT 185.55 35.23 185.71 36.06 ;
      RECT 187.47 37.11 187.63 38.19 ;
      RECT 186.51 36.79 186.67 38.19 ;
      RECT 185.55 37.11 185.71 38.19 ;
      RECT 187.37 36.79 187.53 37.39 ;
      RECT 185.65 36.79 185.81 37.39 ;
      RECT 185.65 36.79 187.53 36.95 ;
      RECT 185.73 68.07 187.55 68.23 ;
      RECT 185.73 62.02 185.89 68.23 ;
      RECT 185.73 62.02 186.11 62.18 ;
      RECT 185.95 57.45 186.11 62.18 ;
      RECT 185.95 57.45 187.55 57.61 ;
      RECT 187.23 57.39 187.55 57.61 ;
      RECT 187.23 53.74 187.39 57.61 ;
      RECT 187.39 51.32 187.55 53.9 ;
      RECT 187.07 51.32 187.55 51.48 ;
      RECT 187.07 49.88 187.23 51.48 ;
      RECT 186.75 49.88 187.23 50.04 ;
      RECT 186.75 47.71 186.91 50.04 ;
      RECT 186.29 47.71 186.91 47.99 ;
      RECT 187.07 47.39 187.23 49.72 ;
      RECT 186.75 47.39 187.23 47.55 ;
      RECT 186.75 43.85 186.91 47.55 ;
      RECT 186.75 43.85 187.53 44.01 ;
      RECT 187.37 39.56 187.53 44.01 ;
      RECT 187.19 39.56 187.53 39.84 ;
      RECT 187.19 39.16 187.35 39.84 ;
      RECT 187.23 62.9 187.39 67.89 ;
      RECT 187.11 64.59 187.39 65.31 ;
      RECT 186.47 52.58 187.23 52.86 ;
      RECT 187.07 51.64 187.23 52.86 ;
      RECT 186.47 52.18 186.63 52.86 ;
      RECT 186.87 34.44 187.21 34.72 ;
      RECT 186.87 32.44 187.03 34.72 ;
      RECT 186.87 33.11 187.21 33.39 ;
      RECT 186.87 32.44 187.21 32.72 ;
      RECT 186.87 40.7 187.21 40.98 ;
      RECT 186.87 38.7 187.03 40.98 ;
      RECT 186.87 40.03 187.21 40.31 ;
      RECT 186.87 38.7 187.21 38.98 ;
      RECT 186.93 53.23 187.21 53.51 ;
      RECT 186.93 53.03 187.09 53.51 ;
      RECT 186.11 53.03 187.09 53.19 ;
      RECT 186.11 50.98 186.27 53.19 ;
      RECT 186.07 52.54 186.27 52.82 ;
      RECT 185.73 50.98 186.27 51.14 ;
      RECT 185.73 50.8 185.95 51.14 ;
      RECT 185.63 56.67 185.79 61.86 ;
      RECT 185.63 56.67 187.07 56.83 ;
      RECT 186.91 56 187.07 56.83 ;
      RECT 185.79 54.4 185.95 56.83 ;
      RECT 186.75 50.66 186.91 51.5 ;
      RECT 186.11 50.66 186.91 50.82 ;
      RECT 186.11 50.18 186.27 50.82 ;
      RECT 185.63 50.18 186.27 50.5 ;
      RECT 185.63 47.07 185.79 50.5 ;
      RECT 185.63 47.07 186.11 47.23 ;
      RECT 185.95 45.44 186.11 47.23 ;
      RECT 186.51 55.68 186.67 56.51 ;
      RECT 186.51 55.68 186.91 55.84 ;
      RECT 186.75 53.67 186.91 55.84 ;
      RECT 186.27 53.67 186.91 53.83 ;
      RECT 186.27 53.35 186.55 53.83 ;
      RECT 186.75 62.9 186.91 67.89 ;
      RECT 186.69 65.82 186.91 66.55 ;
      RECT 186.43 51.7 186.81 51.92 ;
      RECT 186.43 50.98 186.59 51.92 ;
      RECT 185.95 47.39 186.11 49.72 ;
      RECT 185.95 47.39 186.43 47.55 ;
      RECT 186.27 43.85 186.43 47.55 ;
      RECT 185.65 43.85 186.43 44.01 ;
      RECT 185.65 39.56 185.81 44.01 ;
      RECT 185.65 39.56 185.99 39.84 ;
      RECT 185.83 39.16 185.99 39.84 ;
      RECT 185.97 34.44 186.31 34.72 ;
      RECT 186.15 32.44 186.31 34.72 ;
      RECT 185.97 33.11 186.31 33.39 ;
      RECT 185.97 32.44 186.31 32.72 ;
      RECT 185.97 40.7 186.31 40.98 ;
      RECT 186.15 38.7 186.31 40.98 ;
      RECT 185.97 40.03 186.31 40.31 ;
      RECT 185.97 38.7 186.31 38.98 ;
      RECT 186.11 54.06 186.27 56.51 ;
      RECT 185.75 54.06 186.27 54.22 ;
      RECT 185.75 52.98 185.95 54.22 ;
      RECT 185.75 51.34 185.91 54.22 ;
      RECT 185.75 51.34 185.95 52.12 ;
      RECT 185.31 46.75 185.47 47.43 ;
      RECT 184.99 46.75 185.79 46.91 ;
      RECT 185.63 44.23 185.79 46.91 ;
      RECT 184.99 44.23 185.15 46.91 ;
      RECT 183.09 34.88 185.29 35.04 ;
      RECT 185.01 34.59 185.29 35.04 ;
      RECT 184.07 34.59 184.31 35.04 ;
      RECT 183.09 34.59 183.37 35.04 ;
      RECT 184.07 38.38 184.31 39.02 ;
      RECT 185.01 38.38 185.29 38.83 ;
      RECT 183.09 38.38 183.37 38.83 ;
      RECT 183.09 38.38 185.29 38.54 ;
      RECT 183.25 36.47 185.13 36.63 ;
      RECT 184.97 35.86 185.13 36.63 ;
      RECT 184.11 35.23 184.27 36.63 ;
      RECT 183.25 35.86 183.41 36.63 ;
      RECT 185.07 35.23 185.23 36.05 ;
      RECT 183.15 35.23 183.31 36.05 ;
      RECT 185.07 37.11 185.23 38.19 ;
      RECT 184.11 36.79 184.27 38.19 ;
      RECT 183.15 37.11 183.31 38.19 ;
      RECT 184.97 36.79 185.13 37.39 ;
      RECT 183.25 36.79 183.41 37.39 ;
      RECT 183.25 36.79 185.13 36.95 ;
      RECT 183.87 50.66 184.03 51.5 ;
      RECT 183.87 50.66 184.67 50.82 ;
      RECT 184.51 50.18 184.67 50.82 ;
      RECT 184.51 50.18 185.15 50.5 ;
      RECT 184.99 47.07 185.15 50.5 ;
      RECT 184.67 47.07 185.15 47.23 ;
      RECT 184.67 45.44 184.83 47.23 ;
      RECT 184.99 56.67 185.15 61.86 ;
      RECT 183.71 56.67 185.15 56.83 ;
      RECT 184.83 54.4 184.99 56.83 ;
      RECT 183.71 56 183.87 56.83 ;
      RECT 184.67 47.39 184.83 49.72 ;
      RECT 184.35 47.39 184.83 47.55 ;
      RECT 184.35 43.85 184.51 47.55 ;
      RECT 184.35 43.85 185.13 44.01 ;
      RECT 184.97 39.56 185.13 44.01 ;
      RECT 184.79 39.56 185.13 39.84 ;
      RECT 184.79 39.16 184.95 39.84 ;
      RECT 183.57 53.23 183.85 53.51 ;
      RECT 183.69 53.03 183.85 53.51 ;
      RECT 183.69 53.03 184.67 53.19 ;
      RECT 184.51 50.98 184.67 53.19 ;
      RECT 184.51 52.54 184.71 52.82 ;
      RECT 184.51 50.98 185.05 51.14 ;
      RECT 184.83 50.8 185.05 51.14 ;
      RECT 183.23 68.07 185.05 68.23 ;
      RECT 184.89 62.02 185.05 68.23 ;
      RECT 184.67 62.02 185.05 62.18 ;
      RECT 184.67 57.45 184.83 62.18 ;
      RECT 183.23 57.45 184.83 57.61 ;
      RECT 183.23 57.39 183.55 57.61 ;
      RECT 183.39 53.74 183.55 57.61 ;
      RECT 183.23 51.32 183.39 53.9 ;
      RECT 183.23 51.32 183.71 51.48 ;
      RECT 183.55 49.88 183.71 51.48 ;
      RECT 183.55 49.88 184.03 50.04 ;
      RECT 183.87 47.71 184.03 50.04 ;
      RECT 183.87 47.71 184.49 47.99 ;
      RECT 184.51 54.06 184.67 56.51 ;
      RECT 184.51 54.06 185.03 54.22 ;
      RECT 184.87 51.34 185.03 54.22 ;
      RECT 184.83 52.98 185.03 54.22 ;
      RECT 184.83 51.34 185.03 52.12 ;
      RECT 184.47 34.44 184.81 34.72 ;
      RECT 184.47 32.44 184.63 34.72 ;
      RECT 184.47 33.11 184.81 33.39 ;
      RECT 184.47 32.44 184.81 32.72 ;
      RECT 184.47 40.7 184.81 40.98 ;
      RECT 184.47 38.7 184.63 40.98 ;
      RECT 184.47 40.03 184.81 40.31 ;
      RECT 184.47 38.7 184.81 38.98 ;
      RECT 184.11 55.68 184.27 56.51 ;
      RECT 183.87 55.68 184.27 55.84 ;
      RECT 183.87 53.67 184.03 55.84 ;
      RECT 183.87 53.67 184.51 53.83 ;
      RECT 184.23 53.35 184.51 53.83 ;
      RECT 183.97 51.7 184.35 51.92 ;
      RECT 184.19 50.98 184.35 51.92 ;
      RECT 183.55 52.58 184.31 52.86 ;
      RECT 184.15 52.18 184.31 52.86 ;
      RECT 183.55 51.64 183.71 52.86 ;
      RECT 183.87 62.9 184.03 67.89 ;
      RECT 183.87 65.82 184.09 66.55 ;
      RECT 183.55 47.39 183.71 49.72 ;
      RECT 183.55 47.39 184.03 47.55 ;
      RECT 183.87 43.85 184.03 47.55 ;
      RECT 183.25 43.85 184.03 44.01 ;
      RECT 183.25 39.56 183.41 44.01 ;
      RECT 183.25 39.56 183.59 39.84 ;
      RECT 183.43 39.16 183.59 39.84 ;
      RECT 183.57 34.44 183.91 34.72 ;
      RECT 183.75 32.44 183.91 34.72 ;
      RECT 183.57 33.11 183.91 33.39 ;
      RECT 183.57 32.44 183.91 32.72 ;
      RECT 183.57 40.7 183.91 40.98 ;
      RECT 183.75 38.7 183.91 40.98 ;
      RECT 183.57 40.03 183.91 40.31 ;
      RECT 183.57 38.7 183.91 38.98 ;
      RECT 183.39 62.9 183.55 67.89 ;
      RECT 183.39 64.59 183.67 65.31 ;
      RECT 182.91 46.75 183.07 47.43 ;
      RECT 182.59 46.75 183.39 46.91 ;
      RECT 183.23 44.23 183.39 46.91 ;
      RECT 182.59 44.23 182.75 46.91 ;
      RECT 182.39 10.08 182.55 11.89 ;
      RECT 182.39 10.08 183.13 10.24 ;
      RECT 182.91 8.88 183.07 10.24 ;
      RECT 182.91 7.5 183.07 8.72 ;
      RECT 182.86 7.58 183.07 7.9 ;
      RECT 181.83 7.59 183.07 7.75 ;
      RECT 182.79 7.58 183.07 7.75 ;
      RECT 174.87 15.8 175.03 16.08 ;
      RECT 171.75 15.8 171.91 16.08 ;
      RECT 174.27 15.8 175.03 15.96 ;
      RECT 171.75 15.8 172.51 15.96 ;
      RECT 172.35 14.07 172.51 15.96 ;
      RECT 180.77 14.25 180.93 15.89 ;
      RECT 165.85 14.25 166.01 15.89 ;
      RECT 173.31 12.21 173.47 15.8 ;
      RECT 174.27 14.07 174.43 15.96 ;
      RECT 178.25 14.12 178.43 15.79 ;
      RECT 176.97 14.1 177.13 15.79 ;
      RECT 169.65 14.1 169.81 15.79 ;
      RECT 168.35 14.12 168.53 15.79 ;
      RECT 182.11 14.64 182.27 15.6 ;
      RECT 164.51 14.64 164.67 15.6 ;
      RECT 182.91 12.64 183.07 14.96 ;
      RECT 163.71 12.64 163.87 14.96 ;
      RECT 175.93 14.1 176.09 14.89 ;
      RECT 170.69 14.1 170.85 14.89 ;
      RECT 180.49 14.64 183.07 14.84 ;
      RECT 163.71 14.64 166.29 14.84 ;
      RECT 166.13 12.56 166.29 14.84 ;
      RECT 180.49 14.25 181.94 14.84 ;
      RECT 164.84 14.25 166.29 14.84 ;
      RECT 174.99 14.36 176.09 14.52 ;
      RECT 170.69 14.36 171.79 14.52 ;
      RECT 171.63 14.08 171.79 14.52 ;
      RECT 174.99 14.08 175.15 14.52 ;
      RECT 176.97 14.12 180.65 14.28 ;
      RECT 164.84 14.25 169.81 14.28 ;
      RECT 175.93 14.1 177.45 14.26 ;
      RECT 169.33 14.1 170.85 14.26 ;
      RECT 166.13 14.12 170.85 14.26 ;
      RECT 174.27 14.08 175.15 14.24 ;
      RECT 171.63 14.08 172.51 14.24 ;
      RECT 172.17 14.07 174.61 14.23 ;
      RECT 180.49 12.56 180.65 14.84 ;
      RECT 179.53 12.55 179.69 14.28 ;
      RECT 178.65 13.45 178.81 14.28 ;
      RECT 167.97 13.45 168.13 14.28 ;
      RECT 167.09 12.55 167.25 14.28 ;
      RECT 176.19 12.32 176.35 14.26 ;
      RECT 170.43 12.32 170.59 14.26 ;
      RECT 174.45 13.38 174.61 14.24 ;
      RECT 172.17 13.38 172.33 14.24 ;
      RECT 178.57 12.55 178.73 13.61 ;
      RECT 168.05 12.55 168.21 13.61 ;
      RECT 174.33 13.38 174.61 13.54 ;
      RECT 172.17 13.38 172.45 13.54 ;
      RECT 182.24 17.18 182.4 18.9 ;
      RECT 182.24 17.96 183.07 18.12 ;
      RECT 182.91 17.84 183.07 18.12 ;
      RECT 182.2 17.06 182.36 17.34 ;
      RECT 181.22 19.61 181.38 21.25 ;
      RECT 174.27 20.42 174.43 21.25 ;
      RECT 173.31 16.39 173.47 21.25 ;
      RECT 172.35 20.42 172.51 21.25 ;
      RECT 165.4 19.61 165.56 21.25 ;
      RECT 182 20.89 182.42 21.05 ;
      RECT 180.26 19.61 180.42 21.05 ;
      RECT 166.36 19.61 166.52 21.05 ;
      RECT 164.36 20.89 164.78 21.05 ;
      RECT 164.62 19.61 164.78 21.05 ;
      RECT 179.26 20.21 179.42 20.89 ;
      RECT 177.01 20.43 177.17 20.89 ;
      RECT 169.61 20.43 169.77 20.89 ;
      RECT 167.36 20.21 167.52 20.89 ;
      RECT 182 19.61 182.16 21.05 ;
      RECT 176.55 20.43 177.17 20.59 ;
      RECT 169.61 20.43 170.23 20.59 ;
      RECT 170.07 19.1 170.23 20.59 ;
      RECT 174.35 19.16 174.51 20.58 ;
      RECT 172.27 19.16 172.43 20.58 ;
      RECT 175.59 19.16 175.75 20.49 ;
      RECT 171.03 19.16 171.19 20.49 ;
      RECT 176.55 19.1 176.71 20.59 ;
      RECT 179.26 20.21 180.42 20.37 ;
      RECT 180.22 19.61 180.42 20.37 ;
      RECT 166.36 20.21 167.52 20.37 ;
      RECT 166.36 19.61 166.56 20.37 ;
      RECT 180.22 19.61 181.38 19.81 ;
      RECT 165.4 19.61 166.56 19.81 ;
      RECT 180.05 19.61 182.99 19.77 ;
      RECT 163.79 19.61 166.73 19.77 ;
      RECT 166.57 19.1 166.73 19.77 ;
      RECT 179.09 19.1 179.37 19.73 ;
      RECT 167.41 19.1 167.69 19.73 ;
      RECT 180.05 19.1 180.21 19.77 ;
      RECT 175.59 19.16 176.71 19.37 ;
      RECT 170.07 19.16 171.19 19.37 ;
      RECT 170.07 19.16 176.71 19.32 ;
      RECT 175.7 19.1 180.21 19.26 ;
      RECT 175.23 18.46 175.39 19.32 ;
      RECT 174.27 17.56 174.43 19.32 ;
      RECT 172.35 17.56 172.51 19.32 ;
      RECT 171.39 18.46 171.55 19.32 ;
      RECT 166.57 19.1 171.08 19.26 ;
      RECT 169.94 17.76 170.1 19.26 ;
      RECT 176.68 19.01 178.6 19.26 ;
      RECT 178.42 16.65 178.6 19.26 ;
      RECT 168.18 19.01 170.1 19.26 ;
      RECT 177.48 17.58 177.64 19.26 ;
      RECT 176.68 17.76 176.84 19.26 ;
      RECT 169.14 17.58 169.3 19.26 ;
      RECT 168.18 16.65 168.36 19.26 ;
      RECT 176.15 17.76 176.84 17.92 ;
      RECT 169.94 17.76 170.63 17.92 ;
      RECT 170.47 16.77 170.63 17.92 ;
      RECT 176.15 16.77 176.31 17.92 ;
      RECT 182.68 15.57 182.84 17.28 ;
      RECT 182.08 16.43 182.24 16.71 ;
      RECT 182.08 16.43 182.84 16.59 ;
      RECT 182.62 15.57 182.9 15.73 ;
      RECT 180.69 34.88 182.89 35.04 ;
      RECT 182.61 34.59 182.89 35.04 ;
      RECT 181.67 34.59 181.91 35.04 ;
      RECT 180.69 34.59 180.97 35.04 ;
      RECT 181.67 38.38 181.91 39.02 ;
      RECT 182.61 38.38 182.89 38.83 ;
      RECT 180.69 38.38 180.97 38.83 ;
      RECT 180.69 38.38 182.89 38.54 ;
      RECT 182.21 23.66 182.75 23.82 ;
      RECT 182.59 20.12 182.75 23.82 ;
      RECT 182.29 23.22 182.75 23.38 ;
      RECT 182.59 20.83 182.84 21.11 ;
      RECT 182.32 20.12 182.75 20.28 ;
      RECT 182.64 26.15 182.8 28.96 ;
      RECT 182.64 26.15 182.83 26.51 ;
      RECT 180.85 36.47 182.73 36.63 ;
      RECT 182.57 35.88 182.73 36.63 ;
      RECT 181.71 35.23 181.87 36.63 ;
      RECT 180.85 35.88 181.01 36.63 ;
      RECT 182.67 35.23 182.83 36.06 ;
      RECT 180.75 35.23 180.91 36.06 ;
      RECT 182.67 37.11 182.83 38.19 ;
      RECT 181.71 36.79 181.87 38.19 ;
      RECT 180.75 37.11 180.91 38.19 ;
      RECT 182.57 36.79 182.73 37.39 ;
      RECT 180.85 36.79 181.01 37.39 ;
      RECT 180.85 36.79 182.73 36.95 ;
      RECT 180.93 68.07 182.75 68.23 ;
      RECT 180.93 62.02 181.09 68.23 ;
      RECT 180.93 62.02 181.31 62.18 ;
      RECT 181.15 57.45 181.31 62.18 ;
      RECT 181.15 57.45 182.75 57.61 ;
      RECT 182.43 57.39 182.75 57.61 ;
      RECT 182.43 53.74 182.59 57.61 ;
      RECT 182.59 51.32 182.75 53.9 ;
      RECT 182.27 51.32 182.75 51.48 ;
      RECT 182.27 49.88 182.43 51.48 ;
      RECT 181.95 49.88 182.43 50.04 ;
      RECT 181.95 47.71 182.11 50.04 ;
      RECT 181.49 47.71 182.11 47.99 ;
      RECT 182.27 47.39 182.43 49.72 ;
      RECT 181.95 47.39 182.43 47.55 ;
      RECT 181.95 43.85 182.11 47.55 ;
      RECT 181.95 43.85 182.73 44.01 ;
      RECT 182.57 39.56 182.73 44.01 ;
      RECT 182.39 39.56 182.73 39.84 ;
      RECT 182.39 39.16 182.55 39.84 ;
      RECT 180.09 8.96 180.41 9.12 ;
      RECT 180.09 7.8 180.25 9.12 ;
      RECT 182.43 7.91 182.59 8.8 ;
      RECT 181.51 7.91 182.59 8.07 ;
      RECT 180.09 7.8 181.67 7.96 ;
      RECT 182.41 23.98 182.59 24.52 ;
      RECT 181.89 23.98 182.59 24.14 ;
      RECT 181.89 23.27 182.05 24.14 ;
      RECT 181.95 21.78 182.11 23.43 ;
      RECT 181.81 21.21 181.97 21.94 ;
      RECT 181.68 20.95 181.84 21.37 ;
      RECT 182.43 62.9 182.59 67.89 ;
      RECT 182.31 64.59 182.59 65.31 ;
      RECT 181.67 52.58 182.43 52.86 ;
      RECT 182.27 51.64 182.43 52.86 ;
      RECT 181.67 52.18 181.83 52.86 ;
      RECT 182.07 34.44 182.41 34.72 ;
      RECT 182.07 32.44 182.23 34.72 ;
      RECT 182.07 33.11 182.41 33.39 ;
      RECT 182.07 32.44 182.41 32.72 ;
      RECT 182.07 40.7 182.41 40.98 ;
      RECT 182.07 38.7 182.23 40.98 ;
      RECT 182.07 40.03 182.41 40.31 ;
      RECT 182.07 38.7 182.41 38.98 ;
      RECT 182.13 53.23 182.41 53.51 ;
      RECT 182.13 53.03 182.29 53.51 ;
      RECT 181.31 53.03 182.29 53.19 ;
      RECT 181.31 50.98 181.47 53.19 ;
      RECT 181.27 52.54 181.47 52.82 ;
      RECT 180.93 50.98 181.47 51.14 ;
      RECT 180.93 50.8 181.15 51.14 ;
      RECT 181.31 28.52 182.4 28.68 ;
      RECT 181.31 28.35 181.59 28.68 ;
      RECT 180.91 28.35 181.59 28.51 ;
      RECT 182.16 24.79 182.32 28.32 ;
      RECT 181.63 25.16 182.32 25.32 ;
      RECT 182.11 12.92 182.27 13.67 ;
      RECT 181.91 12.92 182.27 13.08 ;
      RECT 181.91 9.68 182.07 13.08 ;
      RECT 181.91 9.68 182.11 11.89 ;
      RECT 181.13 9.68 182.11 9.84 ;
      RECT 181.13 8.6 181.29 9.84 ;
      RECT 180.83 56.67 180.99 61.86 ;
      RECT 180.83 56.67 182.27 56.83 ;
      RECT 182.11 56 182.27 56.83 ;
      RECT 180.99 54.4 181.15 56.83 ;
      RECT 180.27 26.02 180.83 26.18 ;
      RECT 180.67 25.58 180.83 26.18 ;
      RECT 180.67 25.58 181.37 25.74 ;
      RECT 181.21 22.71 181.37 25.74 ;
      RECT 181.17 24 181.37 25.74 ;
      RECT 181.17 24.3 182.17 24.46 ;
      RECT 181.11 22.04 181.27 22.99 ;
      RECT 180.95 21.85 181.11 22.32 ;
      RECT 181.95 50.66 182.11 51.5 ;
      RECT 181.31 50.66 182.11 50.82 ;
      RECT 181.31 50.18 181.47 50.82 ;
      RECT 180.83 50.18 181.47 50.5 ;
      RECT 180.83 47.07 180.99 50.5 ;
      RECT 180.83 47.07 181.31 47.23 ;
      RECT 181.15 45.44 181.31 47.23 ;
      RECT 181.71 55.68 181.87 56.51 ;
      RECT 181.71 55.68 182.11 55.84 ;
      RECT 181.95 53.67 182.11 55.84 ;
      RECT 181.47 53.67 182.11 53.83 ;
      RECT 181.47 53.35 181.75 53.83 ;
      RECT 181.95 62.9 182.11 67.89 ;
      RECT 181.89 65.82 182.11 66.55 ;
      RECT 181.63 51.7 182.01 51.92 ;
      RECT 181.63 50.98 181.79 51.92 ;
      RECT 179.05 26.36 179.21 26.72 ;
      RECT 179.05 26.36 181.35 26.52 ;
      RECT 181.19 26.04 181.35 26.52 ;
      RECT 181.19 26.04 182 26.2 ;
      RECT 181.76 16.52 181.92 18.9 ;
      RECT 181.56 16.52 181.92 16.8 ;
      RECT 181.63 15.31 181.79 16.8 ;
      RECT 181.43 22.13 181.79 22.41 ;
      RECT 181.43 21.53 181.59 22.41 ;
      RECT 180.56 21.53 180.72 21.92 ;
      RECT 180.56 21.53 181.59 21.69 ;
      RECT 180.74 20.21 180.9 21.69 ;
      RECT 181.59 11.5 181.75 13.22 ;
      RECT 180.23 12.22 181.75 12.38 ;
      RECT 181.33 11.5 181.75 11.66 ;
      RECT 181.15 47.39 181.31 49.72 ;
      RECT 181.15 47.39 181.63 47.55 ;
      RECT 181.47 43.85 181.63 47.55 ;
      RECT 180.85 43.85 181.63 44.01 ;
      RECT 180.85 39.56 181.01 44.01 ;
      RECT 180.85 39.56 181.19 39.84 ;
      RECT 181.03 39.16 181.19 39.84 ;
      RECT 180.66 18.3 181.6 18.46 ;
      RECT 181.24 17.05 181.6 18.46 ;
      RECT 181.24 16.2 181.4 18.46 ;
      RECT 180.49 16.2 181.45 16.36 ;
      RECT 181.29 16.08 181.45 16.36 ;
      RECT 180.05 16.07 180.72 16.23 ;
      RECT 181.17 34.44 181.51 34.72 ;
      RECT 181.35 32.44 181.51 34.72 ;
      RECT 181.17 33.11 181.51 33.39 ;
      RECT 181.17 32.44 181.51 32.72 ;
      RECT 181.17 40.7 181.51 40.98 ;
      RECT 181.35 38.7 181.51 40.98 ;
      RECT 181.17 40.03 181.51 40.31 ;
      RECT 181.17 38.7 181.51 38.98 ;
      RECT 181.31 54.06 181.47 56.51 ;
      RECT 180.95 54.06 181.47 54.22 ;
      RECT 180.95 52.98 181.15 54.22 ;
      RECT 180.95 51.34 181.11 54.22 ;
      RECT 180.95 51.34 181.15 52.12 ;
      RECT 179.22 28.01 181.38 28.17 ;
      RECT 181.22 26.68 181.38 28.17 ;
      RECT 180.22 26.97 180.38 28.17 ;
      RECT 179.22 27.93 179.54 28.17 ;
      RECT 179.22 27.34 179.38 28.17 ;
      RECT 180.01 12.56 180.17 13.61 ;
      RECT 179.91 11.9 180.07 13.24 ;
      RECT 179.91 11.9 181.19 12.06 ;
      RECT 180.09 9.6 180.25 12.06 ;
      RECT 180.9 16.52 181.08 16.84 ;
      RECT 180.18 16.52 181.08 16.68 ;
      RECT 180.89 23.18 181.05 23.84 ;
      RECT 180.72 23.18 181.05 23.34 ;
      RECT 180.72 22.65 180.88 23.34 ;
      RECT 180.51 46.75 180.67 47.43 ;
      RECT 180.19 46.75 180.99 46.91 ;
      RECT 180.83 44.23 180.99 46.91 ;
      RECT 180.19 44.23 180.35 46.91 ;
      RECT 180.7 26.69 180.86 27.85 ;
      RECT 180.66 26.69 180.9 27.33 ;
      RECT 180.57 9.28 180.73 11.72 ;
      RECT 179.61 8.12 179.77 11.72 ;
      RECT 178.65 8.5 178.81 11.72 ;
      RECT 176.99 9.63 177.15 11.4 ;
      RECT 176.99 9.95 178.81 10.11 ;
      RECT 177.68 9.79 177.84 10.11 ;
      RECT 180.61 8.12 180.81 9.84 ;
      RECT 176.93 9.63 177.44 9.79 ;
      RECT 179.61 9.28 180.81 9.44 ;
      RECT 178.61 8.5 178.92 8.78 ;
      RECT 178.61 8.56 179.77 8.72 ;
      RECT 175.63 28.74 180.75 28.9 ;
      RECT 178.83 27.92 178.99 28.9 ;
      RECT 177.39 27.92 177.55 28.9 ;
      RECT 180.44 16.92 180.6 18.12 ;
      RECT 180.2 16.92 180.6 17.08 ;
      RECT 178.29 34.88 180.49 35.04 ;
      RECT 180.21 34.59 180.49 35.04 ;
      RECT 179.27 34.59 179.51 35.04 ;
      RECT 178.29 34.59 178.57 35.04 ;
      RECT 179.27 38.38 179.51 39.02 ;
      RECT 180.21 38.38 180.49 38.83 ;
      RECT 178.29 38.38 178.57 38.83 ;
      RECT 178.29 38.38 180.49 38.54 ;
      RECT 178.11 21.69 178.27 26.21 ;
      RECT 179.35 24.34 179.51 26.2 ;
      RECT 176.87 24.35 177.03 26.2 ;
      RECT 180.23 24.04 180.45 25.52 ;
      RECT 175.93 24.04 176.15 25.52 ;
      RECT 179.35 24.46 180.45 24.63 ;
      RECT 175.93 24.46 177.03 24.63 ;
      RECT 176.85 21.69 177.01 24.63 ;
      RECT 179.37 21.69 179.53 24.63 ;
      RECT 176.85 21.69 179.53 21.85 ;
      RECT 178.45 36.47 180.33 36.63 ;
      RECT 180.17 35.86 180.33 36.63 ;
      RECT 179.31 35.23 179.47 36.63 ;
      RECT 178.45 35.86 178.61 36.63 ;
      RECT 180.27 35.23 180.43 36.05 ;
      RECT 178.35 35.23 178.51 36.05 ;
      RECT 180.27 37.11 180.43 38.19 ;
      RECT 179.31 36.79 179.47 38.19 ;
      RECT 178.35 37.11 178.51 38.19 ;
      RECT 180.17 36.79 180.33 37.39 ;
      RECT 178.45 36.79 178.61 37.39 ;
      RECT 178.45 36.79 180.33 36.95 ;
      RECT 180.23 21.37 180.39 23.37 ;
      RECT 176.39 21.37 180.39 21.53 ;
      RECT 179.74 20.73 179.9 21.53 ;
      RECT 176.39 20.78 176.55 21.53 ;
      RECT 179.07 50.66 179.23 51.5 ;
      RECT 179.07 50.66 179.87 50.82 ;
      RECT 179.71 50.18 179.87 50.82 ;
      RECT 179.71 50.18 180.35 50.5 ;
      RECT 180.19 47.07 180.35 50.5 ;
      RECT 179.87 47.07 180.35 47.23 ;
      RECT 179.87 45.44 180.03 47.23 ;
      RECT 180.19 56.67 180.35 61.86 ;
      RECT 178.91 56.67 180.35 56.83 ;
      RECT 180.03 54.4 180.19 56.83 ;
      RECT 178.91 56 179.07 56.83 ;
      RECT 179.87 47.39 180.03 49.72 ;
      RECT 179.55 47.39 180.03 47.55 ;
      RECT 179.55 43.85 179.71 47.55 ;
      RECT 179.55 43.85 180.33 44.01 ;
      RECT 180.17 39.56 180.33 44.01 ;
      RECT 179.99 39.56 180.33 39.84 ;
      RECT 179.99 39.16 180.15 39.84 ;
      RECT 178.77 53.23 179.05 53.51 ;
      RECT 178.89 53.03 179.05 53.51 ;
      RECT 178.89 53.03 179.87 53.19 ;
      RECT 179.71 50.98 179.87 53.19 ;
      RECT 179.71 52.54 179.91 52.82 ;
      RECT 179.71 50.98 180.25 51.14 ;
      RECT 180.03 50.8 180.25 51.14 ;
      RECT 178.43 68.07 180.25 68.23 ;
      RECT 180.09 62.02 180.25 68.23 ;
      RECT 179.87 62.02 180.25 62.18 ;
      RECT 179.87 57.45 180.03 62.18 ;
      RECT 178.43 57.45 180.03 57.61 ;
      RECT 178.43 57.39 178.75 57.61 ;
      RECT 178.59 53.74 178.75 57.61 ;
      RECT 178.43 51.32 178.59 53.9 ;
      RECT 178.43 51.32 178.91 51.48 ;
      RECT 178.75 49.88 178.91 51.48 ;
      RECT 178.75 49.88 179.23 50.04 ;
      RECT 179.07 47.71 179.23 50.04 ;
      RECT 179.07 47.71 179.69 47.99 ;
      RECT 179.71 54.06 179.87 56.51 ;
      RECT 179.71 54.06 180.23 54.22 ;
      RECT 180.07 51.34 180.23 54.22 ;
      RECT 180.03 52.98 180.23 54.22 ;
      RECT 180.03 51.34 180.23 52.12 ;
      RECT 178.92 18.78 180.04 18.94 ;
      RECT 179.86 17.48 180.04 18.94 ;
      RECT 177.96 17.26 178.13 18.8 ;
      RECT 177.97 16.12 178.13 18.8 ;
      RECT 177 16.44 177.16 18.8 ;
      RECT 178.92 16.03 179.08 18.94 ;
      RECT 176.95 16.44 177.16 17.57 ;
      RECT 179.86 16.44 180.02 18.94 ;
      RECT 176.95 17.26 178.13 17.42 ;
      RECT 176.95 16.44 177.23 17.42 ;
      RECT 179.73 14.52 179.89 16.71 ;
      RECT 175.95 16.12 179.08 16.28 ;
      RECT 178.77 14.52 178.93 16.28 ;
      RECT 177.77 14.84 177.93 16.28 ;
      RECT 178.77 14.52 179.89 14.68 ;
      RECT 179.67 34.44 180.01 34.72 ;
      RECT 179.67 32.44 179.83 34.72 ;
      RECT 179.67 33.11 180.01 33.39 ;
      RECT 179.67 32.44 180.01 32.72 ;
      RECT 179.67 40.7 180.01 40.98 ;
      RECT 179.67 38.7 179.83 40.98 ;
      RECT 179.67 40.03 180.01 40.31 ;
      RECT 179.67 38.7 180.01 38.98 ;
      RECT 179.83 21.85 179.99 24.3 ;
      RECT 179.69 21.85 179.99 22.13 ;
      RECT 179.67 24.79 179.87 25.35 ;
      RECT 179.67 24.79 179.99 25.03 ;
      RECT 178.35 28.04 178.67 28.32 ;
      RECT 178.51 25.99 178.67 28.32 ;
      RECT 179.7 27.02 179.86 27.7 ;
      RECT 178.51 27.02 179.86 27.18 ;
      RECT 178.51 25.99 178.89 26.23 ;
      RECT 178.73 25.16 178.89 26.23 ;
      RECT 178.37 20.26 178.53 21.05 ;
      RECT 178.37 20.26 179.1 20.44 ;
      RECT 178.94 19.89 179.1 20.44 ;
      RECT 178.94 19.89 179.76 20.05 ;
      RECT 179.57 19.61 179.76 20.05 ;
      RECT 179.57 19.61 179.85 19.77 ;
      RECT 179.31 55.68 179.47 56.51 ;
      RECT 179.07 55.68 179.47 55.84 ;
      RECT 179.07 53.67 179.23 55.84 ;
      RECT 179.07 53.67 179.71 53.83 ;
      RECT 179.43 53.35 179.71 53.83 ;
      RECT 179.17 51.7 179.55 51.92 ;
      RECT 179.39 50.98 179.55 51.92 ;
      RECT 178.75 52.58 179.51 52.86 ;
      RECT 179.35 52.18 179.51 52.86 ;
      RECT 178.75 51.64 178.91 52.86 ;
      RECT 179.05 12.53 179.21 13.61 ;
      RECT 179.21 11.88 179.37 12.69 ;
      RECT 178.25 11.77 178.49 12.05 ;
      RECT 178.25 11.88 179.37 12.04 ;
      RECT 179.13 8.88 179.29 12.04 ;
      RECT 179.07 62.9 179.23 67.89 ;
      RECT 179.07 65.82 179.29 66.55 ;
      RECT 178.75 47.39 178.91 49.72 ;
      RECT 178.75 47.39 179.23 47.55 ;
      RECT 179.07 43.85 179.23 47.55 ;
      RECT 178.45 43.85 179.23 44.01 ;
      RECT 178.45 39.56 178.61 44.01 ;
      RECT 178.45 39.56 178.79 39.84 ;
      RECT 178.63 39.16 178.79 39.84 ;
      RECT 179.05 22.01 179.21 23.37 ;
      RECT 178.43 22.01 179.21 22.17 ;
      RECT 178.73 24.72 179.11 24.96 ;
      RECT 178.73 22.35 178.89 24.96 ;
      RECT 178.77 34.44 179.11 34.72 ;
      RECT 178.95 32.44 179.11 34.72 ;
      RECT 178.77 33.11 179.11 33.39 ;
      RECT 178.77 32.44 179.11 32.72 ;
      RECT 178.77 40.7 179.11 40.98 ;
      RECT 178.95 38.7 179.11 40.98 ;
      RECT 178.77 40.03 179.11 40.31 ;
      RECT 178.77 38.7 179.11 38.98 ;
      RECT 177.47 12.21 177.63 13.28 ;
      RECT 177.47 12.21 179.05 12.37 ;
      RECT 177.93 11.47 178.09 12.37 ;
      RECT 177.99 10.85 178.15 11.63 ;
      RECT 178.59 62.9 178.75 67.89 ;
      RECT 178.59 64.59 178.87 65.31 ;
      RECT 178.11 46.75 178.27 47.43 ;
      RECT 177.79 46.75 178.59 46.91 ;
      RECT 178.43 44.23 178.59 46.91 ;
      RECT 177.79 44.23 177.95 46.91 ;
      RECT 178.31 10.51 178.47 11.24 ;
      RECT 177.81 10.51 178.47 10.67 ;
      RECT 178.16 8.96 178.32 9.79 ;
      RECT 177.13 8.96 178.32 9.12 ;
      RECT 177.83 20.63 178.11 20.79 ;
      RECT 177.95 19.59 178.11 20.79 ;
      RECT 175.89 34.88 178.09 35.04 ;
      RECT 177.81 34.59 178.09 35.04 ;
      RECT 176.87 34.59 177.11 35.04 ;
      RECT 175.89 34.59 176.17 35.04 ;
      RECT 176.87 38.38 177.11 39.02 ;
      RECT 177.81 38.38 178.09 38.83 ;
      RECT 175.89 38.38 176.17 38.83 ;
      RECT 175.89 38.38 178.09 38.54 ;
      RECT 177.71 28.04 178.03 28.32 ;
      RECT 177.71 25.99 177.87 28.32 ;
      RECT 176.52 27.02 176.68 27.7 ;
      RECT 176.52 27.02 177.87 27.18 ;
      RECT 177.49 25.99 177.87 26.23 ;
      RECT 177.49 25.16 177.65 26.23 ;
      RECT 176.05 36.47 177.93 36.63 ;
      RECT 177.77 35.88 177.93 36.63 ;
      RECT 176.91 35.23 177.07 36.63 ;
      RECT 176.05 35.88 176.21 36.63 ;
      RECT 177.87 35.23 178.03 36.06 ;
      RECT 175.95 35.23 176.11 36.06 ;
      RECT 177.87 37.11 178.03 38.19 ;
      RECT 176.91 36.79 177.07 38.19 ;
      RECT 175.95 37.11 176.11 38.19 ;
      RECT 177.77 36.79 177.93 37.39 ;
      RECT 176.05 36.79 176.21 37.39 ;
      RECT 176.05 36.79 177.93 36.95 ;
      RECT 177.17 22.01 177.33 23.37 ;
      RECT 177.17 22.01 177.95 22.17 ;
      RECT 176.13 68.07 177.95 68.23 ;
      RECT 176.13 62.02 176.29 68.23 ;
      RECT 176.13 62.02 176.51 62.18 ;
      RECT 176.35 57.45 176.51 62.18 ;
      RECT 176.35 57.45 177.95 57.61 ;
      RECT 177.63 57.39 177.95 57.61 ;
      RECT 177.63 53.74 177.79 57.61 ;
      RECT 177.79 51.32 177.95 53.9 ;
      RECT 177.47 51.32 177.95 51.48 ;
      RECT 177.47 49.88 177.63 51.48 ;
      RECT 177.15 49.88 177.63 50.04 ;
      RECT 177.15 47.71 177.31 50.04 ;
      RECT 176.69 47.71 177.31 47.99 ;
      RECT 177.47 47.39 177.63 49.72 ;
      RECT 177.15 47.39 177.63 47.55 ;
      RECT 177.15 43.85 177.31 47.55 ;
      RECT 177.15 43.85 177.93 44.01 ;
      RECT 177.77 39.56 177.93 44.01 ;
      RECT 177.59 39.56 177.93 39.84 ;
      RECT 177.59 39.16 177.75 39.84 ;
      RECT 177.29 14.44 177.45 15.64 ;
      RECT 177.29 14.44 177.79 14.6 ;
      RECT 177.63 62.9 177.79 67.89 ;
      RECT 177.51 64.59 177.79 65.31 ;
      RECT 177.27 24.72 177.65 24.96 ;
      RECT 177.49 22.35 177.65 24.96 ;
      RECT 176.99 12.32 177.15 13.37 ;
      RECT 177.11 11.56 177.27 12.48 ;
      RECT 176.51 11.56 177.63 11.72 ;
      RECT 177.47 10.27 177.63 11.72 ;
      RECT 176.51 10.4 176.67 11.72 ;
      RECT 176.87 52.58 177.63 52.86 ;
      RECT 177.47 51.64 177.63 52.86 ;
      RECT 176.87 52.18 177.03 52.86 ;
      RECT 177.27 34.44 177.61 34.72 ;
      RECT 177.27 32.44 177.43 34.72 ;
      RECT 177.27 33.11 177.61 33.39 ;
      RECT 177.27 32.44 177.61 32.72 ;
      RECT 177.27 40.7 177.61 40.98 ;
      RECT 177.27 38.7 177.43 40.98 ;
      RECT 177.27 40.03 177.61 40.31 ;
      RECT 177.27 38.7 177.61 38.98 ;
      RECT 177.33 53.23 177.61 53.51 ;
      RECT 177.33 53.03 177.49 53.51 ;
      RECT 176.51 53.03 177.49 53.19 ;
      RECT 176.51 50.98 176.67 53.19 ;
      RECT 176.47 52.54 176.67 52.82 ;
      RECT 176.13 50.98 176.67 51.14 ;
      RECT 176.13 50.8 176.35 51.14 ;
      RECT 176.03 56.67 176.19 61.86 ;
      RECT 176.03 56.67 177.47 56.83 ;
      RECT 177.31 56 177.47 56.83 ;
      RECT 176.19 54.4 176.35 56.83 ;
      RECT 177.17 26.36 177.33 26.72 ;
      RECT 175.03 26.36 177.33 26.52 ;
      RECT 175.03 26.04 175.19 26.52 ;
      RECT 174.38 26.04 175.19 26.2 ;
      RECT 177.15 50.66 177.31 51.5 ;
      RECT 176.51 50.66 177.31 50.82 ;
      RECT 176.51 50.18 176.67 50.82 ;
      RECT 176.03 50.18 176.67 50.5 ;
      RECT 176.03 47.07 176.19 50.5 ;
      RECT 176.03 47.07 176.51 47.23 ;
      RECT 176.35 45.44 176.51 47.23 ;
      RECT 176.91 55.68 177.07 56.51 ;
      RECT 176.91 55.68 177.31 55.84 ;
      RECT 177.15 53.67 177.31 55.84 ;
      RECT 176.67 53.67 177.31 53.83 ;
      RECT 176.67 53.35 176.95 53.83 ;
      RECT 177.15 62.9 177.31 67.89 ;
      RECT 177.09 65.82 177.31 66.55 ;
      RECT 176.83 51.7 177.21 51.92 ;
      RECT 176.83 50.98 176.99 51.92 ;
      RECT 175 28.01 177.16 28.17 ;
      RECT 177 27.34 177.16 28.17 ;
      RECT 176.84 27.93 177.16 28.17 ;
      RECT 176 26.97 176.16 28.17 ;
      RECT 175 26.68 175.16 28.17 ;
      RECT 176.51 12 176.67 12.84 ;
      RECT 176.51 12 176.95 12.16 ;
      RECT 176.79 11.88 176.95 12.16 ;
      RECT 175.26 8.82 176.85 8.98 ;
      RECT 176.69 7.16 176.85 8.98 ;
      RECT 176.35 47.39 176.51 49.72 ;
      RECT 176.35 47.39 176.83 47.55 ;
      RECT 176.67 43.85 176.83 47.55 ;
      RECT 176.05 43.85 176.83 44.01 ;
      RECT 176.05 39.56 176.21 44.01 ;
      RECT 176.05 39.56 176.39 39.84 ;
      RECT 176.23 39.16 176.39 39.84 ;
      RECT 176.66 9.92 176.82 10.24 ;
      RECT 176.42 9.92 176.82 10.12 ;
      RECT 175.63 15.8 175.79 17.77 ;
      RECT 175.63 15.8 176.45 15.96 ;
      RECT 176.45 14.42 176.61 15.88 ;
      RECT 176.27 15.72 176.61 15.88 ;
      RECT 176.45 14.42 176.79 14.58 ;
      RECT 176.51 24.79 176.71 25.35 ;
      RECT 176.39 24.79 176.71 25.03 ;
      RECT 176.37 34.44 176.71 34.72 ;
      RECT 176.55 32.44 176.71 34.72 ;
      RECT 176.37 33.11 176.71 33.39 ;
      RECT 176.37 32.44 176.71 32.72 ;
      RECT 176.37 40.7 176.71 40.98 ;
      RECT 176.55 38.7 176.71 40.98 ;
      RECT 176.37 40.03 176.71 40.31 ;
      RECT 176.37 38.7 176.71 38.98 ;
      RECT 176.39 21.85 176.55 24.3 ;
      RECT 176.39 21.85 176.69 22.13 ;
      RECT 176.51 54.06 176.67 56.51 ;
      RECT 176.15 54.06 176.67 54.22 ;
      RECT 176.15 52.98 176.35 54.22 ;
      RECT 176.15 51.34 176.31 54.22 ;
      RECT 176.15 51.34 176.35 52.12 ;
      RECT 176.01 18.51 176.2 18.94 ;
      RECT 175.81 18.51 176.5 18.7 ;
      RECT 175.99 21.29 176.15 23.37 ;
      RECT 176.07 19.81 176.23 21.46 ;
      RECT 175.61 12.58 175.89 13.24 ;
      RECT 175.73 11.84 175.89 13.24 ;
      RECT 175.37 11.84 175.53 12.12 ;
      RECT 175.37 11.84 176.21 12 ;
      RECT 176.05 10.46 176.21 12 ;
      RECT 175.71 46.75 175.87 47.43 ;
      RECT 175.39 46.75 176.19 46.91 ;
      RECT 176.03 44.23 176.19 46.91 ;
      RECT 175.39 44.23 175.55 46.91 ;
      RECT 175.55 26.02 176.11 26.18 ;
      RECT 175.55 25.58 175.71 26.18 ;
      RECT 175.01 25.58 175.71 25.74 ;
      RECT 175.01 24 175.21 25.74 ;
      RECT 174.27 24.24 175.21 24.52 ;
      RECT 174.27 21.85 174.43 24.52 ;
      RECT 174.94 9.14 175.13 9.52 ;
      RECT 174.94 9.14 176.07 9.3 ;
      RECT 174.94 8.52 175.1 9.52 ;
      RECT 174.92 8.36 175.08 8.64 ;
      RECT 175.31 18.13 175.97 18.3 ;
      RECT 175.31 15 175.47 18.3 ;
      RECT 175.31 15.32 176.01 15.64 ;
      RECT 174.85 15 175.47 15.16 ;
      RECT 175.57 9.68 175.73 11.68 ;
      RECT 171.05 9.68 171.21 11.68 ;
      RECT 174.11 9.68 174.27 11.36 ;
      RECT 172.51 9.68 172.67 11.36 ;
      RECT 172.51 10.76 174.27 10.92 ;
      RECT 173.31 8.38 173.47 10.92 ;
      RECT 174.11 9.68 175.73 9.84 ;
      RECT 175.45 9.46 175.61 9.84 ;
      RECT 171.05 9.68 172.67 9.84 ;
      RECT 171.17 9.46 171.33 9.84 ;
      RECT 175.52 26.68 175.68 27.85 ;
      RECT 175.48 26.68 175.72 27.33 ;
      RECT 173.49 34.88 175.69 35.04 ;
      RECT 175.41 34.59 175.69 35.04 ;
      RECT 174.47 34.59 174.71 35.04 ;
      RECT 173.49 34.59 173.77 35.04 ;
      RECT 174.47 38.38 174.71 39.02 ;
      RECT 175.41 38.38 175.69 38.83 ;
      RECT 173.49 38.38 173.77 38.83 ;
      RECT 173.49 38.38 175.69 38.54 ;
      RECT 175.47 13.5 175.63 14.2 ;
      RECT 175.29 13.5 175.63 13.66 ;
      RECT 175.29 12.52 175.45 13.66 ;
      RECT 175.05 12.52 175.45 12.84 ;
      RECT 175.05 10.84 175.21 12.84 ;
      RECT 173.65 36.47 175.53 36.63 ;
      RECT 175.37 35.86 175.53 36.63 ;
      RECT 174.51 35.23 174.67 36.63 ;
      RECT 173.65 35.86 173.81 36.63 ;
      RECT 175.47 35.23 175.63 36.05 ;
      RECT 173.55 35.23 173.71 36.05 ;
      RECT 175.47 37.11 175.63 38.19 ;
      RECT 174.51 36.79 174.67 38.19 ;
      RECT 173.55 37.11 173.71 38.19 ;
      RECT 175.37 36.79 175.53 37.39 ;
      RECT 173.65 36.79 173.81 37.39 ;
      RECT 173.65 36.79 175.53 36.95 ;
      RECT 174.27 50.66 174.43 51.5 ;
      RECT 174.27 50.66 175.07 50.82 ;
      RECT 174.91 50.18 175.07 50.82 ;
      RECT 174.91 50.18 175.55 50.5 ;
      RECT 175.39 47.07 175.55 50.5 ;
      RECT 175.07 47.07 175.55 47.23 ;
      RECT 175.07 45.44 175.23 47.23 ;
      RECT 175.39 56.67 175.55 61.86 ;
      RECT 174.11 56.67 175.55 56.83 ;
      RECT 175.23 54.4 175.39 56.83 ;
      RECT 174.11 56 174.27 56.83 ;
      RECT 175.07 47.39 175.23 49.72 ;
      RECT 174.75 47.39 175.23 47.55 ;
      RECT 174.75 43.85 174.91 47.55 ;
      RECT 174.75 43.85 175.53 44.01 ;
      RECT 175.37 39.56 175.53 44.01 ;
      RECT 175.19 39.56 175.53 39.84 ;
      RECT 175.19 39.16 175.35 39.84 ;
      RECT 175.33 23.12 175.49 23.84 ;
      RECT 174.59 23.12 175.49 23.28 ;
      RECT 174.59 20.86 174.75 23.28 ;
      RECT 174.59 20.86 174.95 21.02 ;
      RECT 174.79 20.74 174.95 21.02 ;
      RECT 173.98 28.52 175.07 28.68 ;
      RECT 174.79 28.35 175.07 28.68 ;
      RECT 174.79 28.35 175.47 28.51 ;
      RECT 173.97 53.23 174.25 53.51 ;
      RECT 174.09 53.03 174.25 53.51 ;
      RECT 174.09 53.03 175.07 53.19 ;
      RECT 174.91 50.98 175.07 53.19 ;
      RECT 174.91 52.54 175.11 52.82 ;
      RECT 174.91 50.98 175.45 51.14 ;
      RECT 175.23 50.8 175.45 51.14 ;
      RECT 173.63 68.07 175.45 68.23 ;
      RECT 175.29 62.02 175.45 68.23 ;
      RECT 175.07 62.02 175.45 62.18 ;
      RECT 175.07 57.45 175.23 62.18 ;
      RECT 173.63 57.45 175.23 57.61 ;
      RECT 173.63 57.39 173.95 57.61 ;
      RECT 173.79 53.74 173.95 57.61 ;
      RECT 173.63 51.32 173.79 53.9 ;
      RECT 173.63 51.32 174.11 51.48 ;
      RECT 173.95 49.88 174.11 51.48 ;
      RECT 173.95 49.88 174.43 50.04 ;
      RECT 174.27 47.71 174.43 50.04 ;
      RECT 174.27 47.71 174.89 47.99 ;
      RECT 174.91 54.06 175.07 56.51 ;
      RECT 174.91 54.06 175.43 54.22 ;
      RECT 175.27 51.34 175.43 54.22 ;
      RECT 175.23 52.98 175.43 54.22 ;
      RECT 175.23 51.34 175.43 52.12 ;
      RECT 174.87 13.06 175.03 13.54 ;
      RECT 174.59 13.06 175.03 13.22 ;
      RECT 174.59 10 174.75 13.22 ;
      RECT 174.59 10 175.41 10.16 ;
      RECT 174.95 22.29 175.19 22.53 ;
      RECT 174.95 21.18 175.11 22.53 ;
      RECT 174.91 21.18 175.11 21.58 ;
      RECT 175.11 19.81 175.28 21.35 ;
      RECT 174.87 34.44 175.21 34.72 ;
      RECT 174.87 32.44 175.03 34.72 ;
      RECT 174.87 33.11 175.21 33.39 ;
      RECT 174.87 32.44 175.21 32.72 ;
      RECT 174.87 40.7 175.21 40.98 ;
      RECT 174.87 38.7 175.03 40.98 ;
      RECT 174.87 40.03 175.21 40.31 ;
      RECT 174.87 38.7 175.21 38.98 ;
      RECT 174.75 17.24 174.91 19 ;
      RECT 173.79 14.39 173.95 18.85 ;
      RECT 173.79 17.24 174.91 17.4 ;
      RECT 173.77 15.32 173.97 16.04 ;
      RECT 173.79 14.39 173.97 16.04 ;
      RECT 174.51 55.68 174.67 56.51 ;
      RECT 174.27 55.68 174.67 55.84 ;
      RECT 174.27 53.67 174.43 55.84 ;
      RECT 174.27 53.67 174.91 53.83 ;
      RECT 174.63 53.35 174.91 53.83 ;
      RECT 174.06 24.7 174.22 28.32 ;
      RECT 174.06 25.16 174.75 25.32 ;
      RECT 173.53 24.7 174.22 24.86 ;
      RECT 174.37 51.7 174.75 51.92 ;
      RECT 174.59 50.98 174.75 51.92 ;
      RECT 173.95 52.58 174.71 52.86 ;
      RECT 174.55 52.18 174.71 52.86 ;
      RECT 173.95 51.64 174.11 52.86 ;
      RECT 174.27 62.9 174.43 67.89 ;
      RECT 174.27 65.82 174.49 66.55 ;
      RECT 173.71 9.36 173.87 10.6 ;
      RECT 173.71 9.36 174.45 9.52 ;
      RECT 173.95 47.39 174.11 49.72 ;
      RECT 173.95 47.39 174.43 47.55 ;
      RECT 174.27 43.85 174.43 47.55 ;
      RECT 173.65 43.85 174.43 44.01 ;
      RECT 173.65 39.56 173.81 44.01 ;
      RECT 173.65 39.56 173.99 39.84 ;
      RECT 173.83 39.16 173.99 39.84 ;
      RECT 173.97 34.44 174.31 34.72 ;
      RECT 174.15 32.44 174.31 34.72 ;
      RECT 173.97 33.11 174.31 33.39 ;
      RECT 173.97 32.44 174.31 32.72 ;
      RECT 173.97 40.7 174.31 40.98 ;
      RECT 174.15 38.7 174.31 40.98 ;
      RECT 173.97 40.03 174.31 40.31 ;
      RECT 173.97 38.7 174.31 38.98 ;
      RECT 173.87 11.52 174.03 12.43 ;
      RECT 173.87 11.75 174.11 12.03 ;
      RECT 173.59 11.52 174.03 11.68 ;
      RECT 173.59 11.08 173.75 11.68 ;
      RECT 173.79 62.9 173.95 67.89 ;
      RECT 173.79 64.59 174.07 65.31 ;
      RECT 173.79 23.73 173.97 24.54 ;
      RECT 173.79 20.48 173.95 24.54 ;
      RECT 173.31 46.75 173.47 47.43 ;
      RECT 172.99 46.75 173.79 46.91 ;
      RECT 173.63 44.23 173.79 46.91 ;
      RECT 172.99 44.23 173.15 46.91 ;
      RECT 173.58 26.15 173.74 28.96 ;
      RECT 173.55 26.15 173.74 26.51 ;
      RECT 171.09 34.88 173.29 35.04 ;
      RECT 173.01 34.59 173.29 35.04 ;
      RECT 172.07 34.59 172.31 35.04 ;
      RECT 171.09 34.59 171.37 35.04 ;
      RECT 172.07 38.38 172.31 39.02 ;
      RECT 173.01 38.38 173.29 38.83 ;
      RECT 171.09 38.38 171.37 38.83 ;
      RECT 171.09 38.38 173.29 38.54 ;
      RECT 172.56 24.7 172.72 28.32 ;
      RECT 172.03 25.16 172.72 25.32 ;
      RECT 172.56 24.7 173.25 24.86 ;
      RECT 173.04 26.15 173.2 28.96 ;
      RECT 173.04 26.15 173.23 26.51 ;
      RECT 171.25 36.47 173.13 36.63 ;
      RECT 172.97 35.88 173.13 36.63 ;
      RECT 172.11 35.23 172.27 36.63 ;
      RECT 171.25 35.88 171.41 36.63 ;
      RECT 173.07 35.23 173.23 36.06 ;
      RECT 171.15 35.23 171.31 36.06 ;
      RECT 173.07 37.11 173.23 38.19 ;
      RECT 172.11 36.79 172.27 38.19 ;
      RECT 171.15 37.11 171.31 38.19 ;
      RECT 172.97 36.79 173.13 37.39 ;
      RECT 171.25 36.79 171.41 37.39 ;
      RECT 171.25 36.79 173.13 36.95 ;
      RECT 172.75 11.52 172.91 12.43 ;
      RECT 172.67 11.75 172.91 12.03 ;
      RECT 172.75 11.52 173.19 11.68 ;
      RECT 173.03 11.08 173.19 11.68 ;
      RECT 171.33 68.07 173.15 68.23 ;
      RECT 171.33 62.02 171.49 68.23 ;
      RECT 171.33 62.02 171.71 62.18 ;
      RECT 171.55 57.45 171.71 62.18 ;
      RECT 171.55 57.45 173.15 57.61 ;
      RECT 172.83 57.39 173.15 57.61 ;
      RECT 172.83 53.74 172.99 57.61 ;
      RECT 172.99 51.32 173.15 53.9 ;
      RECT 172.67 51.32 173.15 51.48 ;
      RECT 172.67 49.88 172.83 51.48 ;
      RECT 172.35 49.88 172.83 50.04 ;
      RECT 172.35 47.71 172.51 50.04 ;
      RECT 171.89 47.71 172.51 47.99 ;
      RECT 172.67 47.39 172.83 49.72 ;
      RECT 172.35 47.39 172.83 47.55 ;
      RECT 172.35 43.85 172.51 47.55 ;
      RECT 172.35 43.85 173.13 44.01 ;
      RECT 172.97 39.56 173.13 44.01 ;
      RECT 172.79 39.56 173.13 39.84 ;
      RECT 172.79 39.16 172.95 39.84 ;
      RECT 172.91 9.36 173.07 10.6 ;
      RECT 172.33 9.36 173.07 9.52 ;
      RECT 171.87 17.24 172.03 19 ;
      RECT 172.83 14.39 172.99 18.85 ;
      RECT 171.87 17.24 172.99 17.4 ;
      RECT 172.81 15.32 173.01 16.04 ;
      RECT 172.81 14.39 172.99 16.04 ;
      RECT 172.81 23.73 172.99 24.54 ;
      RECT 172.83 20.48 172.99 24.54 ;
      RECT 172.83 62.9 172.99 67.89 ;
      RECT 172.71 64.59 172.99 65.31 ;
      RECT 172.07 52.58 172.83 52.86 ;
      RECT 172.67 51.64 172.83 52.86 ;
      RECT 172.07 52.18 172.23 52.86 ;
      RECT 172.47 34.44 172.81 34.72 ;
      RECT 172.47 32.44 172.63 34.72 ;
      RECT 172.47 33.11 172.81 33.39 ;
      RECT 172.47 32.44 172.81 32.72 ;
      RECT 172.47 40.7 172.81 40.98 ;
      RECT 172.47 38.7 172.63 40.98 ;
      RECT 172.47 40.03 172.81 40.31 ;
      RECT 172.47 38.7 172.81 38.98 ;
      RECT 172.53 53.23 172.81 53.51 ;
      RECT 172.53 53.03 172.69 53.51 ;
      RECT 171.71 53.03 172.69 53.19 ;
      RECT 171.71 50.98 171.87 53.19 ;
      RECT 171.67 52.54 171.87 52.82 ;
      RECT 171.33 50.98 171.87 51.14 ;
      RECT 171.33 50.8 171.55 51.14 ;
      RECT 171.71 28.52 172.8 28.68 ;
      RECT 171.71 28.35 171.99 28.68 ;
      RECT 171.31 28.35 171.99 28.51 ;
      RECT 171.23 56.67 171.39 61.86 ;
      RECT 171.23 56.67 172.67 56.83 ;
      RECT 172.51 56 172.67 56.83 ;
      RECT 171.39 54.4 171.55 56.83 ;
      RECT 170.67 26.02 171.23 26.18 ;
      RECT 171.07 25.58 171.23 26.18 ;
      RECT 171.07 25.58 171.77 25.74 ;
      RECT 171.57 24 171.77 25.74 ;
      RECT 171.57 24.24 172.51 24.52 ;
      RECT 172.35 21.85 172.51 24.52 ;
      RECT 172.35 50.66 172.51 51.5 ;
      RECT 171.71 50.66 172.51 50.82 ;
      RECT 171.71 50.18 171.87 50.82 ;
      RECT 171.23 50.18 171.87 50.5 ;
      RECT 171.23 47.07 171.39 50.5 ;
      RECT 171.23 47.07 171.71 47.23 ;
      RECT 171.55 45.44 171.71 47.23 ;
      RECT 172.11 55.68 172.27 56.51 ;
      RECT 172.11 55.68 172.51 55.84 ;
      RECT 172.35 53.67 172.51 55.84 ;
      RECT 171.87 53.67 172.51 53.83 ;
      RECT 171.87 53.35 172.15 53.83 ;
      RECT 172.35 62.9 172.51 67.89 ;
      RECT 172.29 65.82 172.51 66.55 ;
      RECT 172.03 51.7 172.41 51.92 ;
      RECT 172.03 50.98 172.19 51.92 ;
      RECT 169.45 26.36 169.61 26.72 ;
      RECT 169.45 26.36 171.75 26.52 ;
      RECT 171.59 26.04 171.75 26.52 ;
      RECT 171.59 26.04 172.4 26.2 ;
      RECT 171.75 13.06 171.91 13.54 ;
      RECT 171.75 13.06 172.19 13.22 ;
      RECT 172.03 10 172.19 13.22 ;
      RECT 171.37 10 172.19 10.16 ;
      RECT 171.29 23.12 171.45 23.84 ;
      RECT 171.29 23.12 172.19 23.28 ;
      RECT 172.03 20.86 172.19 23.28 ;
      RECT 171.83 20.86 172.19 21.02 ;
      RECT 171.83 20.74 171.99 21.02 ;
      RECT 171.55 47.39 171.71 49.72 ;
      RECT 171.55 47.39 172.03 47.55 ;
      RECT 171.87 43.85 172.03 47.55 ;
      RECT 171.25 43.85 172.03 44.01 ;
      RECT 171.25 39.56 171.41 44.01 ;
      RECT 171.25 39.56 171.59 39.84 ;
      RECT 171.43 39.16 171.59 39.84 ;
      RECT 170.81 18.13 171.47 18.3 ;
      RECT 171.31 15 171.47 18.3 ;
      RECT 170.77 15.32 171.47 15.64 ;
      RECT 171.31 15 171.93 15.16 ;
      RECT 171.57 34.44 171.91 34.72 ;
      RECT 171.75 32.44 171.91 34.72 ;
      RECT 171.57 33.11 171.91 33.39 ;
      RECT 171.57 32.44 171.91 32.72 ;
      RECT 171.57 40.7 171.91 40.98 ;
      RECT 171.75 38.7 171.91 40.98 ;
      RECT 171.57 40.03 171.91 40.31 ;
      RECT 171.57 38.7 171.91 38.98 ;
      RECT 171.59 22.29 171.83 22.53 ;
      RECT 171.67 21.18 171.83 22.53 ;
      RECT 171.67 21.18 171.87 21.58 ;
      RECT 171.5 19.81 171.67 21.35 ;
      RECT 171.71 54.06 171.87 56.51 ;
      RECT 171.35 54.06 171.87 54.22 ;
      RECT 171.35 52.98 171.55 54.22 ;
      RECT 171.35 51.34 171.51 54.22 ;
      RECT 171.35 51.34 171.55 52.12 ;
      RECT 171.65 9.14 171.84 9.52 ;
      RECT 170.71 9.14 171.84 9.3 ;
      RECT 171.68 8.52 171.84 9.52 ;
      RECT 171.7 8.36 171.86 8.64 ;
      RECT 169.62 28.01 171.78 28.17 ;
      RECT 171.62 26.68 171.78 28.17 ;
      RECT 170.62 26.97 170.78 28.17 ;
      RECT 169.62 27.93 169.94 28.17 ;
      RECT 169.62 27.34 169.78 28.17 ;
      RECT 171.15 13.5 171.31 14.2 ;
      RECT 171.15 13.5 171.49 13.66 ;
      RECT 171.33 12.52 171.49 13.66 ;
      RECT 171.33 12.52 171.73 12.84 ;
      RECT 171.57 10.84 171.73 12.84 ;
      RECT 169.93 8.82 171.52 8.98 ;
      RECT 169.93 7.16 170.09 8.98 ;
      RECT 170.89 12.58 171.17 13.24 ;
      RECT 170.89 11.84 171.05 13.24 ;
      RECT 171.25 11.84 171.41 12.12 ;
      RECT 170.57 11.84 171.41 12 ;
      RECT 170.57 10.46 170.73 12 ;
      RECT 170.91 46.75 171.07 47.43 ;
      RECT 170.59 46.75 171.39 46.91 ;
      RECT 171.23 44.23 171.39 46.91 ;
      RECT 170.59 44.23 170.75 46.91 ;
      RECT 171.1 26.68 171.26 27.85 ;
      RECT 171.06 26.68 171.3 27.33 ;
      RECT 170.99 15.8 171.15 17.77 ;
      RECT 170.33 15.8 171.15 15.96 ;
      RECT 170.17 14.42 170.33 15.88 ;
      RECT 170.17 15.72 170.51 15.88 ;
      RECT 169.99 14.42 170.33 14.58 ;
      RECT 166.03 28.74 171.15 28.9 ;
      RECT 169.23 27.92 169.39 28.9 ;
      RECT 167.79 27.92 167.95 28.9 ;
      RECT 170.58 18.51 170.77 18.94 ;
      RECT 170.28 18.51 170.97 18.7 ;
      RECT 168.69 34.88 170.89 35.04 ;
      RECT 170.61 34.59 170.89 35.04 ;
      RECT 169.67 34.59 169.91 35.04 ;
      RECT 168.69 34.59 168.97 35.04 ;
      RECT 169.67 38.38 169.91 39.02 ;
      RECT 170.61 38.38 170.89 38.83 ;
      RECT 168.69 38.38 168.97 38.83 ;
      RECT 168.69 38.38 170.89 38.54 ;
      RECT 168.51 21.69 168.67 26.21 ;
      RECT 169.75 24.35 169.91 26.2 ;
      RECT 167.27 24.34 167.43 26.2 ;
      RECT 170.63 24.04 170.85 25.52 ;
      RECT 166.33 24.04 166.55 25.52 ;
      RECT 169.75 24.46 170.85 24.63 ;
      RECT 166.33 24.46 167.43 24.63 ;
      RECT 167.25 21.69 167.41 24.63 ;
      RECT 169.77 21.69 169.93 24.63 ;
      RECT 167.25 21.69 169.93 21.85 ;
      RECT 166.74 18.78 167.86 18.94 ;
      RECT 169.62 16.44 169.78 18.8 ;
      RECT 168.65 17.26 168.82 18.8 ;
      RECT 167.7 16.03 167.86 18.94 ;
      RECT 166.74 17.48 166.92 18.94 ;
      RECT 169.62 16.44 169.83 17.57 ;
      RECT 166.76 16.44 166.92 18.94 ;
      RECT 168.65 17.26 169.83 17.42 ;
      RECT 169.55 16.44 169.83 17.42 ;
      RECT 168.65 16.12 168.81 18.8 ;
      RECT 166.89 14.52 167.05 16.71 ;
      RECT 167.7 16.12 170.83 16.28 ;
      RECT 168.85 14.84 169.01 16.28 ;
      RECT 167.85 14.52 168.01 16.28 ;
      RECT 166.89 14.52 168.01 14.68 ;
      RECT 168.85 36.47 170.73 36.63 ;
      RECT 170.57 35.86 170.73 36.63 ;
      RECT 169.71 35.23 169.87 36.63 ;
      RECT 168.85 35.86 169.01 36.63 ;
      RECT 170.67 35.23 170.83 36.05 ;
      RECT 168.75 35.23 168.91 36.05 ;
      RECT 170.67 37.11 170.83 38.19 ;
      RECT 169.71 36.79 169.87 38.19 ;
      RECT 168.75 37.11 168.91 38.19 ;
      RECT 170.57 36.79 170.73 37.39 ;
      RECT 168.85 36.79 169.01 37.39 ;
      RECT 168.85 36.79 170.73 36.95 ;
      RECT 170.63 21.29 170.79 23.37 ;
      RECT 170.55 19.81 170.71 21.46 ;
      RECT 169.47 50.66 169.63 51.5 ;
      RECT 169.47 50.66 170.27 50.82 ;
      RECT 170.11 50.18 170.27 50.82 ;
      RECT 170.11 50.18 170.75 50.5 ;
      RECT 170.59 47.07 170.75 50.5 ;
      RECT 170.27 47.07 170.75 47.23 ;
      RECT 170.27 45.44 170.43 47.23 ;
      RECT 170.59 56.67 170.75 61.86 ;
      RECT 169.31 56.67 170.75 56.83 ;
      RECT 170.43 54.4 170.59 56.83 ;
      RECT 169.31 56 169.47 56.83 ;
      RECT 170.27 47.39 170.43 49.72 ;
      RECT 169.95 47.39 170.43 47.55 ;
      RECT 169.95 43.85 170.11 47.55 ;
      RECT 169.95 43.85 170.73 44.01 ;
      RECT 170.57 39.56 170.73 44.01 ;
      RECT 170.39 39.56 170.73 39.84 ;
      RECT 170.39 39.16 170.55 39.84 ;
      RECT 169.17 53.23 169.45 53.51 ;
      RECT 169.29 53.03 169.45 53.51 ;
      RECT 169.29 53.03 170.27 53.19 ;
      RECT 170.11 50.98 170.27 53.19 ;
      RECT 170.11 52.54 170.31 52.82 ;
      RECT 170.11 50.98 170.65 51.14 ;
      RECT 170.43 50.8 170.65 51.14 ;
      RECT 168.83 68.07 170.65 68.23 ;
      RECT 170.49 62.02 170.65 68.23 ;
      RECT 170.27 62.02 170.65 62.18 ;
      RECT 170.27 57.45 170.43 62.18 ;
      RECT 168.83 57.45 170.43 57.61 ;
      RECT 168.83 57.39 169.15 57.61 ;
      RECT 168.99 53.74 169.15 57.61 ;
      RECT 168.83 51.32 168.99 53.9 ;
      RECT 168.83 51.32 169.31 51.48 ;
      RECT 169.15 49.88 169.31 51.48 ;
      RECT 169.15 49.88 169.63 50.04 ;
      RECT 169.47 47.71 169.63 50.04 ;
      RECT 169.47 47.71 170.09 47.99 ;
      RECT 170.11 54.06 170.27 56.51 ;
      RECT 170.11 54.06 170.63 54.22 ;
      RECT 170.47 51.34 170.63 54.22 ;
      RECT 170.43 52.98 170.63 54.22 ;
      RECT 170.43 51.34 170.63 52.12 ;
      RECT 170.07 34.44 170.41 34.72 ;
      RECT 170.07 32.44 170.23 34.72 ;
      RECT 170.07 33.11 170.41 33.39 ;
      RECT 170.07 32.44 170.41 32.72 ;
      RECT 170.07 40.7 170.41 40.98 ;
      RECT 170.07 38.7 170.23 40.98 ;
      RECT 170.07 40.03 170.41 40.31 ;
      RECT 170.07 38.7 170.41 38.98 ;
      RECT 166.39 21.37 166.55 23.37 ;
      RECT 166.39 21.37 170.39 21.53 ;
      RECT 170.23 20.78 170.39 21.53 ;
      RECT 166.88 20.73 167.04 21.53 ;
      RECT 170.23 21.85 170.39 24.3 ;
      RECT 170.09 21.85 170.39 22.13 ;
      RECT 170.07 24.79 170.27 25.35 ;
      RECT 170.07 24.79 170.39 25.03 ;
      RECT 169.96 9.92 170.12 10.24 ;
      RECT 169.96 9.92 170.36 10.12 ;
      RECT 169.63 12.32 169.79 13.37 ;
      RECT 169.51 11.56 169.67 12.48 ;
      RECT 169.15 11.56 170.27 11.72 ;
      RECT 170.11 10.4 170.27 11.72 ;
      RECT 169.15 10.27 169.31 11.72 ;
      RECT 170.11 12 170.27 12.84 ;
      RECT 169.83 12 170.27 12.16 ;
      RECT 169.83 11.88 169.99 12.16 ;
      RECT 168.75 28.04 169.07 28.32 ;
      RECT 168.91 25.99 169.07 28.32 ;
      RECT 170.1 27.02 170.26 27.7 ;
      RECT 168.91 27.02 170.26 27.18 ;
      RECT 168.91 25.99 169.29 26.23 ;
      RECT 169.13 25.16 169.29 26.23 ;
      RECT 169.71 55.68 169.87 56.51 ;
      RECT 169.47 55.68 169.87 55.84 ;
      RECT 169.47 53.67 169.63 55.84 ;
      RECT 169.47 53.67 170.11 53.83 ;
      RECT 169.83 53.35 170.11 53.83 ;
      RECT 169.57 51.7 169.95 51.92 ;
      RECT 169.79 50.98 169.95 51.92 ;
      RECT 169.15 52.58 169.91 52.86 ;
      RECT 169.75 52.18 169.91 52.86 ;
      RECT 169.15 51.64 169.31 52.86 ;
      RECT 167.97 8.5 168.13 11.72 ;
      RECT 167.01 8.12 167.17 11.72 ;
      RECT 166.05 9.28 166.21 11.72 ;
      RECT 169.63 9.63 169.79 11.4 ;
      RECT 167.97 9.95 169.79 10.11 ;
      RECT 168.94 9.79 169.1 10.11 ;
      RECT 165.97 8.12 166.17 9.84 ;
      RECT 169.34 9.63 169.85 9.79 ;
      RECT 165.97 9.28 167.17 9.44 ;
      RECT 167.86 8.5 168.17 8.78 ;
      RECT 167.01 8.56 168.17 8.72 ;
      RECT 169.47 62.9 169.63 67.89 ;
      RECT 169.47 65.82 169.69 66.55 ;
      RECT 168.46 8.96 168.62 9.79 ;
      RECT 168.46 8.96 169.65 9.12 ;
      RECT 169.15 47.39 169.31 49.72 ;
      RECT 169.15 47.39 169.63 47.55 ;
      RECT 169.47 43.85 169.63 47.55 ;
      RECT 168.85 43.85 169.63 44.01 ;
      RECT 168.85 39.56 169.01 44.01 ;
      RECT 168.85 39.56 169.19 39.84 ;
      RECT 169.03 39.16 169.19 39.84 ;
      RECT 169.45 22.01 169.61 23.37 ;
      RECT 168.83 22.01 169.61 22.17 ;
      RECT 169.13 24.72 169.51 24.96 ;
      RECT 169.13 22.35 169.29 24.96 ;
      RECT 169.17 34.44 169.51 34.72 ;
      RECT 169.35 32.44 169.51 34.72 ;
      RECT 169.17 33.11 169.51 33.39 ;
      RECT 169.17 32.44 169.51 32.72 ;
      RECT 169.17 40.7 169.51 40.98 ;
      RECT 169.35 38.7 169.51 40.98 ;
      RECT 169.17 40.03 169.51 40.31 ;
      RECT 169.17 38.7 169.51 38.98 ;
      RECT 169.33 14.44 169.49 15.64 ;
      RECT 168.99 14.44 169.49 14.6 ;
      RECT 169.15 12.21 169.31 13.28 ;
      RECT 167.73 12.21 169.31 12.37 ;
      RECT 168.69 11.47 168.85 12.37 ;
      RECT 168.63 10.85 168.79 11.63 ;
      RECT 168.99 62.9 169.15 67.89 ;
      RECT 168.99 64.59 169.27 65.31 ;
      RECT 168.51 46.75 168.67 47.43 ;
      RECT 168.19 46.75 168.99 46.91 ;
      RECT 168.83 44.23 168.99 46.91 ;
      RECT 168.19 44.23 168.35 46.91 ;
      RECT 168.31 10.51 168.47 11.24 ;
      RECT 168.31 10.51 168.97 10.67 ;
      RECT 168.67 20.63 168.95 20.79 ;
      RECT 168.67 19.59 168.83 20.79 ;
      RECT 167.57 12.53 167.73 13.61 ;
      RECT 167.41 11.88 167.57 12.69 ;
      RECT 168.29 11.77 168.53 12.05 ;
      RECT 167.41 11.88 168.53 12.04 ;
      RECT 167.49 8.88 167.65 12.04 ;
      RECT 166.29 34.88 168.49 35.04 ;
      RECT 168.21 34.59 168.49 35.04 ;
      RECT 167.27 34.59 167.51 35.04 ;
      RECT 166.29 34.59 166.57 35.04 ;
      RECT 167.27 38.38 167.51 39.02 ;
      RECT 168.21 38.38 168.49 38.83 ;
      RECT 166.29 38.38 166.57 38.83 ;
      RECT 166.29 38.38 168.49 38.54 ;
      RECT 168.11 28.04 168.43 28.32 ;
      RECT 168.11 25.99 168.27 28.32 ;
      RECT 166.92 27.02 167.08 27.7 ;
      RECT 166.92 27.02 168.27 27.18 ;
      RECT 167.89 25.99 168.27 26.23 ;
      RECT 167.89 25.16 168.05 26.23 ;
      RECT 166.45 36.47 168.33 36.63 ;
      RECT 168.17 35.88 168.33 36.63 ;
      RECT 167.31 35.23 167.47 36.63 ;
      RECT 166.45 35.88 166.61 36.63 ;
      RECT 168.27 35.23 168.43 36.06 ;
      RECT 166.35 35.23 166.51 36.06 ;
      RECT 168.27 37.11 168.43 38.19 ;
      RECT 167.31 36.79 167.47 38.19 ;
      RECT 166.35 37.11 166.51 38.19 ;
      RECT 168.17 36.79 168.33 37.39 ;
      RECT 166.45 36.79 166.61 37.39 ;
      RECT 166.45 36.79 168.33 36.95 ;
      RECT 168.25 20.26 168.41 21.05 ;
      RECT 167.68 20.26 168.41 20.44 ;
      RECT 167.68 19.89 167.84 20.44 ;
      RECT 167.02 19.89 167.84 20.05 ;
      RECT 167.02 19.61 167.21 20.05 ;
      RECT 166.93 19.61 167.21 19.77 ;
      RECT 167.57 22.01 167.73 23.37 ;
      RECT 167.57 22.01 168.35 22.17 ;
      RECT 166.53 68.07 168.35 68.23 ;
      RECT 166.53 62.02 166.69 68.23 ;
      RECT 166.53 62.02 166.91 62.18 ;
      RECT 166.75 57.45 166.91 62.18 ;
      RECT 166.75 57.45 168.35 57.61 ;
      RECT 168.03 57.39 168.35 57.61 ;
      RECT 168.03 53.74 168.19 57.61 ;
      RECT 168.19 51.32 168.35 53.9 ;
      RECT 167.87 51.32 168.35 51.48 ;
      RECT 167.87 49.88 168.03 51.48 ;
      RECT 167.55 49.88 168.03 50.04 ;
      RECT 167.55 47.71 167.71 50.04 ;
      RECT 167.09 47.71 167.71 47.99 ;
      RECT 167.87 47.39 168.03 49.72 ;
      RECT 167.55 47.39 168.03 47.55 ;
      RECT 167.55 43.85 167.71 47.55 ;
      RECT 167.55 43.85 168.33 44.01 ;
      RECT 168.17 39.56 168.33 44.01 ;
      RECT 167.99 39.56 168.33 39.84 ;
      RECT 167.99 39.16 168.15 39.84 ;
      RECT 168.03 62.9 168.19 67.89 ;
      RECT 167.91 64.59 168.19 65.31 ;
      RECT 167.67 24.72 168.05 24.96 ;
      RECT 167.89 22.35 168.05 24.96 ;
      RECT 167.27 52.58 168.03 52.86 ;
      RECT 167.87 51.64 168.03 52.86 ;
      RECT 167.27 52.18 167.43 52.86 ;
      RECT 167.67 34.44 168.01 34.72 ;
      RECT 167.67 32.44 167.83 34.72 ;
      RECT 167.67 33.11 168.01 33.39 ;
      RECT 167.67 32.44 168.01 32.72 ;
      RECT 167.67 40.7 168.01 40.98 ;
      RECT 167.67 38.7 167.83 40.98 ;
      RECT 167.67 40.03 168.01 40.31 ;
      RECT 167.67 38.7 168.01 38.98 ;
      RECT 167.73 53.23 168.01 53.51 ;
      RECT 167.73 53.03 167.89 53.51 ;
      RECT 166.91 53.03 167.89 53.19 ;
      RECT 166.91 50.98 167.07 53.19 ;
      RECT 166.87 52.54 167.07 52.82 ;
      RECT 166.53 50.98 167.07 51.14 ;
      RECT 166.53 50.8 166.75 51.14 ;
      RECT 166.43 56.67 166.59 61.86 ;
      RECT 166.43 56.67 167.87 56.83 ;
      RECT 167.71 56 167.87 56.83 ;
      RECT 166.59 54.4 166.75 56.83 ;
      RECT 167.57 26.36 167.73 26.72 ;
      RECT 165.43 26.36 167.73 26.52 ;
      RECT 165.43 26.04 165.59 26.52 ;
      RECT 164.78 26.04 165.59 26.2 ;
      RECT 167.55 50.66 167.71 51.5 ;
      RECT 166.91 50.66 167.71 50.82 ;
      RECT 166.91 50.18 167.07 50.82 ;
      RECT 166.43 50.18 167.07 50.5 ;
      RECT 166.43 47.07 166.59 50.5 ;
      RECT 166.43 47.07 166.91 47.23 ;
      RECT 166.75 45.44 166.91 47.23 ;
      RECT 167.31 55.68 167.47 56.51 ;
      RECT 167.31 55.68 167.71 55.84 ;
      RECT 167.55 53.67 167.71 55.84 ;
      RECT 167.07 53.67 167.71 53.83 ;
      RECT 167.07 53.35 167.35 53.83 ;
      RECT 167.55 62.9 167.71 67.89 ;
      RECT 167.49 65.82 167.71 66.55 ;
      RECT 167.23 51.7 167.61 51.92 ;
      RECT 167.23 50.98 167.39 51.92 ;
      RECT 165.4 28.01 167.56 28.17 ;
      RECT 167.4 27.34 167.56 28.17 ;
      RECT 167.24 27.93 167.56 28.17 ;
      RECT 166.4 26.97 166.56 28.17 ;
      RECT 165.4 26.68 165.56 28.17 ;
      RECT 166.75 47.39 166.91 49.72 ;
      RECT 166.75 47.39 167.23 47.55 ;
      RECT 167.07 43.85 167.23 47.55 ;
      RECT 166.45 43.85 167.23 44.01 ;
      RECT 166.45 39.56 166.61 44.01 ;
      RECT 166.45 39.56 166.79 39.84 ;
      RECT 166.63 39.16 166.79 39.84 ;
      RECT 166.91 24.79 167.11 25.35 ;
      RECT 166.79 24.79 167.11 25.03 ;
      RECT 166.77 34.44 167.11 34.72 ;
      RECT 166.95 32.44 167.11 34.72 ;
      RECT 166.77 33.11 167.11 33.39 ;
      RECT 166.77 32.44 167.11 32.72 ;
      RECT 166.77 40.7 167.11 40.98 ;
      RECT 166.95 38.7 167.11 40.98 ;
      RECT 166.77 40.03 167.11 40.31 ;
      RECT 166.77 38.7 167.11 38.98 ;
      RECT 166.79 21.85 166.95 24.3 ;
      RECT 166.79 21.85 167.09 22.13 ;
      RECT 166.91 54.06 167.07 56.51 ;
      RECT 166.55 54.06 167.07 54.22 ;
      RECT 166.55 52.98 166.75 54.22 ;
      RECT 166.55 51.34 166.71 54.22 ;
      RECT 166.55 51.34 166.75 52.12 ;
      RECT 166.61 12.56 166.77 13.61 ;
      RECT 166.71 11.9 166.87 13.24 ;
      RECT 165.59 11.9 166.87 12.06 ;
      RECT 166.53 9.6 166.69 12.06 ;
      RECT 165.18 18.3 166.12 18.46 ;
      RECT 165.18 17.05 165.54 18.46 ;
      RECT 165.38 16.2 165.54 18.46 ;
      RECT 165.33 16.2 166.29 16.36 ;
      RECT 166.06 16.07 166.73 16.23 ;
      RECT 165.33 16.08 165.49 16.36 ;
      RECT 166.37 8.96 166.69 9.12 ;
      RECT 166.53 7.8 166.69 9.12 ;
      RECT 164.19 7.91 164.35 8.8 ;
      RECT 164.19 7.91 165.27 8.07 ;
      RECT 165.11 7.8 166.69 7.96 ;
      RECT 165.7 16.52 165.88 16.84 ;
      RECT 165.7 16.52 166.6 16.68 ;
      RECT 166.11 46.75 166.27 47.43 ;
      RECT 165.79 46.75 166.59 46.91 ;
      RECT 166.43 44.23 166.59 46.91 ;
      RECT 165.79 44.23 165.95 46.91 ;
      RECT 166.18 16.92 166.34 18.12 ;
      RECT 166.18 16.92 166.58 17.08 ;
      RECT 165.03 11.5 165.19 13.22 ;
      RECT 165.03 12.22 166.55 12.38 ;
      RECT 165.03 11.5 165.45 11.66 ;
      RECT 165.95 26.02 166.51 26.18 ;
      RECT 165.95 25.58 166.11 26.18 ;
      RECT 165.41 25.58 166.11 25.74 ;
      RECT 165.41 24 165.61 25.74 ;
      RECT 164.61 24.3 165.61 24.46 ;
      RECT 165.41 22.71 165.57 25.74 ;
      RECT 165.51 22.04 165.67 22.99 ;
      RECT 165.67 21.85 165.83 22.32 ;
      RECT 164.99 22.13 165.35 22.41 ;
      RECT 165.19 21.53 165.35 22.41 ;
      RECT 166.06 21.53 166.22 21.92 ;
      RECT 165.19 21.53 166.22 21.69 ;
      RECT 165.88 20.21 166.04 21.69 ;
      RECT 165.92 26.69 166.08 27.85 ;
      RECT 165.88 26.69 166.12 27.33 ;
      RECT 163.89 34.88 166.09 35.04 ;
      RECT 165.81 34.59 166.09 35.04 ;
      RECT 164.87 34.59 165.11 35.04 ;
      RECT 163.89 34.59 164.17 35.04 ;
      RECT 164.87 38.38 165.11 39.02 ;
      RECT 165.81 38.38 166.09 38.83 ;
      RECT 163.89 38.38 164.17 38.83 ;
      RECT 163.89 38.38 166.09 38.54 ;
      RECT 165.73 23.18 165.89 23.84 ;
      RECT 165.73 23.18 166.06 23.34 ;
      RECT 165.9 22.65 166.06 23.34 ;
      RECT 164.05 36.47 165.93 36.63 ;
      RECT 165.77 35.86 165.93 36.63 ;
      RECT 164.91 35.23 165.07 36.63 ;
      RECT 164.05 35.86 164.21 36.63 ;
      RECT 165.87 35.23 166.03 36.05 ;
      RECT 163.95 35.23 164.11 36.05 ;
      RECT 165.87 37.11 166.03 38.19 ;
      RECT 164.91 36.79 165.07 38.19 ;
      RECT 163.95 37.11 164.11 38.19 ;
      RECT 165.77 36.79 165.93 37.39 ;
      RECT 164.05 36.79 164.21 37.39 ;
      RECT 164.05 36.79 165.93 36.95 ;
      RECT 164.67 50.66 164.83 51.5 ;
      RECT 164.67 50.66 165.47 50.82 ;
      RECT 165.31 50.18 165.47 50.82 ;
      RECT 165.31 50.18 165.95 50.5 ;
      RECT 165.79 47.07 165.95 50.5 ;
      RECT 165.47 47.07 165.95 47.23 ;
      RECT 165.47 45.44 165.63 47.23 ;
      RECT 165.79 56.67 165.95 61.86 ;
      RECT 164.51 56.67 165.95 56.83 ;
      RECT 165.63 54.4 165.79 56.83 ;
      RECT 164.51 56 164.67 56.83 ;
      RECT 165.47 47.39 165.63 49.72 ;
      RECT 165.15 47.39 165.63 47.55 ;
      RECT 165.15 43.85 165.31 47.55 ;
      RECT 165.15 43.85 165.93 44.01 ;
      RECT 165.77 39.56 165.93 44.01 ;
      RECT 165.59 39.56 165.93 39.84 ;
      RECT 165.59 39.16 165.75 39.84 ;
      RECT 164.38 28.52 165.47 28.68 ;
      RECT 165.19 28.35 165.47 28.68 ;
      RECT 165.19 28.35 165.87 28.51 ;
      RECT 164.37 53.23 164.65 53.51 ;
      RECT 164.49 53.03 164.65 53.51 ;
      RECT 164.49 53.03 165.47 53.19 ;
      RECT 165.31 50.98 165.47 53.19 ;
      RECT 165.31 52.54 165.51 52.82 ;
      RECT 165.31 50.98 165.85 51.14 ;
      RECT 165.63 50.8 165.85 51.14 ;
      RECT 164.03 68.07 165.85 68.23 ;
      RECT 165.69 62.02 165.85 68.23 ;
      RECT 165.47 62.02 165.85 62.18 ;
      RECT 165.47 57.45 165.63 62.18 ;
      RECT 164.03 57.45 165.63 57.61 ;
      RECT 164.03 57.39 164.35 57.61 ;
      RECT 164.19 53.74 164.35 57.61 ;
      RECT 164.03 51.32 164.19 53.9 ;
      RECT 164.03 51.32 164.51 51.48 ;
      RECT 164.35 49.88 164.51 51.48 ;
      RECT 164.35 49.88 164.83 50.04 ;
      RECT 164.67 47.71 164.83 50.04 ;
      RECT 164.67 47.71 165.29 47.99 ;
      RECT 165.31 54.06 165.47 56.51 ;
      RECT 165.31 54.06 165.83 54.22 ;
      RECT 165.67 51.34 165.83 54.22 ;
      RECT 165.63 52.98 165.83 54.22 ;
      RECT 165.63 51.34 165.83 52.12 ;
      RECT 164.51 12.92 164.67 13.67 ;
      RECT 164.51 12.92 164.87 13.08 ;
      RECT 164.71 9.68 164.87 13.08 ;
      RECT 164.67 9.68 164.87 11.89 ;
      RECT 164.67 9.68 165.65 9.84 ;
      RECT 165.49 8.6 165.65 9.84 ;
      RECT 165.27 34.44 165.61 34.72 ;
      RECT 165.27 32.44 165.43 34.72 ;
      RECT 165.27 33.11 165.61 33.39 ;
      RECT 165.27 32.44 165.61 32.72 ;
      RECT 165.27 40.7 165.61 40.98 ;
      RECT 165.27 38.7 165.43 40.98 ;
      RECT 165.27 40.03 165.61 40.31 ;
      RECT 165.27 38.7 165.61 38.98 ;
      RECT 164.91 55.68 165.07 56.51 ;
      RECT 164.67 55.68 165.07 55.84 ;
      RECT 164.67 53.67 164.83 55.84 ;
      RECT 164.67 53.67 165.31 53.83 ;
      RECT 165.03 53.35 165.31 53.83 ;
      RECT 164.86 16.52 165.02 18.9 ;
      RECT 164.86 16.52 165.22 16.8 ;
      RECT 164.99 15.31 165.15 16.8 ;
      RECT 164.46 24.79 164.62 28.32 ;
      RECT 164.46 25.16 165.15 25.32 ;
      RECT 164.77 51.7 165.15 51.92 ;
      RECT 164.99 50.98 165.15 51.92 ;
      RECT 164.35 52.58 165.11 52.86 ;
      RECT 164.95 52.18 165.11 52.86 ;
      RECT 164.35 51.64 164.51 52.86 ;
      RECT 164.19 23.98 164.37 24.52 ;
      RECT 164.19 23.98 164.89 24.14 ;
      RECT 164.73 23.27 164.89 24.14 ;
      RECT 164.67 21.78 164.83 23.43 ;
      RECT 164.81 21.21 164.97 21.94 ;
      RECT 164.94 20.95 165.1 21.37 ;
      RECT 163.71 7.5 163.87 8.72 ;
      RECT 163.71 7.58 163.92 7.9 ;
      RECT 163.71 7.59 164.95 7.75 ;
      RECT 163.71 7.58 163.99 7.75 ;
      RECT 164.67 62.9 164.83 67.89 ;
      RECT 164.67 65.82 164.89 66.55 ;
      RECT 164.35 47.39 164.51 49.72 ;
      RECT 164.35 47.39 164.83 47.55 ;
      RECT 164.67 43.85 164.83 47.55 ;
      RECT 164.05 43.85 164.83 44.01 ;
      RECT 164.05 39.56 164.21 44.01 ;
      RECT 164.05 39.56 164.39 39.84 ;
      RECT 164.23 39.16 164.39 39.84 ;
      RECT 164.37 34.44 164.71 34.72 ;
      RECT 164.55 32.44 164.71 34.72 ;
      RECT 164.37 33.11 164.71 33.39 ;
      RECT 164.37 32.44 164.71 32.72 ;
      RECT 164.37 40.7 164.71 40.98 ;
      RECT 164.55 38.7 164.71 40.98 ;
      RECT 164.37 40.03 164.71 40.31 ;
      RECT 164.37 38.7 164.71 38.98 ;
      RECT 163.94 15.57 164.1 17.28 ;
      RECT 164.54 16.43 164.7 16.71 ;
      RECT 163.94 16.43 164.7 16.59 ;
      RECT 163.88 15.57 164.16 15.73 ;
      RECT 164.38 17.18 164.54 18.9 ;
      RECT 163.71 17.96 164.54 18.12 ;
      RECT 163.71 17.84 163.87 18.12 ;
      RECT 164.42 17.06 164.58 17.34 ;
      RECT 164.03 23.66 164.57 23.82 ;
      RECT 164.03 20.12 164.19 23.82 ;
      RECT 164.03 23.22 164.49 23.38 ;
      RECT 163.94 20.83 164.19 21.11 ;
      RECT 164.03 20.12 164.46 20.28 ;
      RECT 164.19 62.9 164.35 67.89 ;
      RECT 164.19 64.59 164.47 65.31 ;
      RECT 164.23 10.08 164.39 11.89 ;
      RECT 163.65 10.08 164.39 10.24 ;
      RECT 163.71 8.88 163.87 10.24 ;
      RECT 163.71 46.75 163.87 47.43 ;
      RECT 163.39 46.75 164.19 46.91 ;
      RECT 164.03 44.23 164.19 46.91 ;
      RECT 163.39 44.23 163.55 46.91 ;
      RECT 163.98 26.15 164.14 28.96 ;
      RECT 163.95 26.15 164.14 26.51 ;
      RECT 161.49 34.88 163.69 35.04 ;
      RECT 163.41 34.59 163.69 35.04 ;
      RECT 162.47 34.59 162.71 35.04 ;
      RECT 161.49 34.59 161.77 35.04 ;
      RECT 162.47 38.38 162.71 39.02 ;
      RECT 163.41 38.38 163.69 38.83 ;
      RECT 161.49 38.38 161.77 38.83 ;
      RECT 161.49 38.38 163.69 38.54 ;
      RECT 161.65 36.47 163.53 36.63 ;
      RECT 163.37 35.88 163.53 36.63 ;
      RECT 162.51 35.23 162.67 36.63 ;
      RECT 161.65 35.88 161.81 36.63 ;
      RECT 163.47 35.23 163.63 36.06 ;
      RECT 161.55 35.23 161.71 36.06 ;
      RECT 163.47 37.11 163.63 38.19 ;
      RECT 162.51 36.79 162.67 38.19 ;
      RECT 161.55 37.11 161.71 38.19 ;
      RECT 163.37 36.79 163.53 37.39 ;
      RECT 161.65 36.79 161.81 37.39 ;
      RECT 161.65 36.79 163.53 36.95 ;
      RECT 161.73 68.07 163.55 68.23 ;
      RECT 161.73 62.02 161.89 68.23 ;
      RECT 161.73 62.02 162.11 62.18 ;
      RECT 161.95 57.45 162.11 62.18 ;
      RECT 161.95 57.45 163.55 57.61 ;
      RECT 163.23 57.39 163.55 57.61 ;
      RECT 163.23 53.74 163.39 57.61 ;
      RECT 163.39 51.32 163.55 53.9 ;
      RECT 163.07 51.32 163.55 51.48 ;
      RECT 163.07 49.88 163.23 51.48 ;
      RECT 162.75 49.88 163.23 50.04 ;
      RECT 162.75 47.71 162.91 50.04 ;
      RECT 162.29 47.71 162.91 47.99 ;
      RECT 163.07 47.39 163.23 49.72 ;
      RECT 162.75 47.39 163.23 47.55 ;
      RECT 162.75 43.85 162.91 47.55 ;
      RECT 162.75 43.85 163.53 44.01 ;
      RECT 163.37 39.56 163.53 44.01 ;
      RECT 163.19 39.56 163.53 39.84 ;
      RECT 163.19 39.16 163.35 39.84 ;
      RECT 163.23 62.9 163.39 67.89 ;
      RECT 163.11 64.59 163.39 65.31 ;
      RECT 162.47 52.58 163.23 52.86 ;
      RECT 163.07 51.64 163.23 52.86 ;
      RECT 162.47 52.18 162.63 52.86 ;
      RECT 162.87 34.44 163.21 34.72 ;
      RECT 162.87 32.44 163.03 34.72 ;
      RECT 162.87 33.11 163.21 33.39 ;
      RECT 162.87 32.44 163.21 32.72 ;
      RECT 162.87 40.7 163.21 40.98 ;
      RECT 162.87 38.7 163.03 40.98 ;
      RECT 162.87 40.03 163.21 40.31 ;
      RECT 162.87 38.7 163.21 38.98 ;
      RECT 162.93 53.23 163.21 53.51 ;
      RECT 162.93 53.03 163.09 53.51 ;
      RECT 162.11 53.03 163.09 53.19 ;
      RECT 162.11 50.98 162.27 53.19 ;
      RECT 162.07 52.54 162.27 52.82 ;
      RECT 161.73 50.98 162.27 51.14 ;
      RECT 161.73 50.8 161.95 51.14 ;
      RECT 161.63 56.67 161.79 61.86 ;
      RECT 161.63 56.67 163.07 56.83 ;
      RECT 162.91 56 163.07 56.83 ;
      RECT 161.79 54.4 161.95 56.83 ;
      RECT 155.07 12.95 162.91 13.55 ;
      RECT 162.31 8.34 162.91 13.55 ;
      RECT 155.07 8.34 155.67 13.55 ;
      RECT 155.07 8.34 162.91 8.88 ;
      RECT 155.07 26.87 162.91 27.47 ;
      RECT 162.31 18.71 162.91 27.47 ;
      RECT 155.07 18.71 155.67 27.47 ;
      RECT 155.07 24.41 162.91 25.01 ;
      RECT 155.07 18.71 162.91 19.31 ;
      RECT 162.75 50.66 162.91 51.5 ;
      RECT 162.11 50.66 162.91 50.82 ;
      RECT 162.11 50.18 162.27 50.82 ;
      RECT 161.63 50.18 162.27 50.5 ;
      RECT 161.63 47.07 161.79 50.5 ;
      RECT 161.63 47.07 162.11 47.23 ;
      RECT 161.95 45.44 162.11 47.23 ;
      RECT 162.51 55.68 162.67 56.51 ;
      RECT 162.51 55.68 162.91 55.84 ;
      RECT 162.75 53.67 162.91 55.84 ;
      RECT 162.27 53.67 162.91 53.83 ;
      RECT 162.27 53.35 162.55 53.83 ;
      RECT 162.75 62.9 162.91 67.89 ;
      RECT 162.69 65.82 162.91 66.55 ;
      RECT 162.43 51.7 162.81 51.92 ;
      RECT 162.43 50.98 162.59 51.92 ;
      RECT 161.95 47.39 162.11 49.72 ;
      RECT 161.95 47.39 162.43 47.55 ;
      RECT 162.27 43.85 162.43 47.55 ;
      RECT 161.65 43.85 162.43 44.01 ;
      RECT 161.65 39.56 161.81 44.01 ;
      RECT 161.65 39.56 161.99 39.84 ;
      RECT 161.83 39.16 161.99 39.84 ;
      RECT 161.97 34.44 162.31 34.72 ;
      RECT 162.15 32.44 162.31 34.72 ;
      RECT 161.97 33.11 162.31 33.39 ;
      RECT 161.97 32.44 162.31 32.72 ;
      RECT 161.97 40.7 162.31 40.98 ;
      RECT 162.15 38.7 162.31 40.98 ;
      RECT 161.97 40.03 162.31 40.31 ;
      RECT 161.97 38.7 162.31 38.98 ;
      RECT 162.11 54.06 162.27 56.51 ;
      RECT 161.75 54.06 162.27 54.22 ;
      RECT 161.75 52.98 161.95 54.22 ;
      RECT 161.75 51.34 161.91 54.22 ;
      RECT 161.75 51.34 161.95 52.12 ;
      RECT 161.31 46.75 161.47 47.43 ;
      RECT 160.99 46.75 161.79 46.91 ;
      RECT 161.63 44.23 161.79 46.91 ;
      RECT 160.99 44.23 161.15 46.91 ;
      RECT 159.09 34.88 161.29 35.04 ;
      RECT 161.01 34.59 161.29 35.04 ;
      RECT 160.07 34.59 160.31 35.04 ;
      RECT 159.09 34.59 159.37 35.04 ;
      RECT 160.07 38.38 160.31 39.02 ;
      RECT 161.01 38.38 161.29 38.83 ;
      RECT 159.09 38.38 159.37 38.83 ;
      RECT 159.09 38.38 161.29 38.54 ;
      RECT 159.25 36.47 161.13 36.63 ;
      RECT 160.97 35.86 161.13 36.63 ;
      RECT 160.11 35.23 160.27 36.63 ;
      RECT 159.25 35.86 159.41 36.63 ;
      RECT 161.07 35.23 161.23 36.05 ;
      RECT 159.15 35.23 159.31 36.05 ;
      RECT 161.07 37.11 161.23 38.19 ;
      RECT 160.11 36.79 160.27 38.19 ;
      RECT 159.15 37.11 159.31 38.19 ;
      RECT 160.97 36.79 161.13 37.39 ;
      RECT 159.25 36.79 159.41 37.39 ;
      RECT 159.25 36.79 161.13 36.95 ;
      RECT 159.87 50.66 160.03 51.5 ;
      RECT 159.87 50.66 160.67 50.82 ;
      RECT 160.51 50.18 160.67 50.82 ;
      RECT 160.51 50.18 161.15 50.5 ;
      RECT 160.99 47.07 161.15 50.5 ;
      RECT 160.67 47.07 161.15 47.23 ;
      RECT 160.67 45.44 160.83 47.23 ;
      RECT 160.99 56.67 161.15 61.86 ;
      RECT 159.71 56.67 161.15 56.83 ;
      RECT 160.83 54.4 160.99 56.83 ;
      RECT 159.71 56 159.87 56.83 ;
      RECT 160.67 47.39 160.83 49.72 ;
      RECT 160.35 47.39 160.83 47.55 ;
      RECT 160.35 43.85 160.51 47.55 ;
      RECT 160.35 43.85 161.13 44.01 ;
      RECT 160.97 39.56 161.13 44.01 ;
      RECT 160.79 39.56 161.13 39.84 ;
      RECT 160.79 39.16 160.95 39.84 ;
      RECT 159.57 53.23 159.85 53.51 ;
      RECT 159.69 53.03 159.85 53.51 ;
      RECT 159.69 53.03 160.67 53.19 ;
      RECT 160.51 50.98 160.67 53.19 ;
      RECT 160.51 52.54 160.71 52.82 ;
      RECT 160.51 50.98 161.05 51.14 ;
      RECT 160.83 50.8 161.05 51.14 ;
      RECT 159.23 68.07 161.05 68.23 ;
      RECT 160.89 62.02 161.05 68.23 ;
      RECT 160.67 62.02 161.05 62.18 ;
      RECT 160.67 57.45 160.83 62.18 ;
      RECT 159.23 57.45 160.83 57.61 ;
      RECT 159.23 57.39 159.55 57.61 ;
      RECT 159.39 53.74 159.55 57.61 ;
      RECT 159.23 51.32 159.39 53.9 ;
      RECT 159.23 51.32 159.71 51.48 ;
      RECT 159.55 49.88 159.71 51.48 ;
      RECT 159.55 49.88 160.03 50.04 ;
      RECT 159.87 47.71 160.03 50.04 ;
      RECT 159.87 47.71 160.49 47.99 ;
      RECT 160.51 54.06 160.67 56.51 ;
      RECT 160.51 54.06 161.03 54.22 ;
      RECT 160.87 51.34 161.03 54.22 ;
      RECT 160.83 52.98 161.03 54.22 ;
      RECT 160.83 51.34 161.03 52.12 ;
      RECT 160.47 34.44 160.81 34.72 ;
      RECT 160.47 32.44 160.63 34.72 ;
      RECT 160.47 33.11 160.81 33.39 ;
      RECT 160.47 32.44 160.81 32.72 ;
      RECT 160.47 40.7 160.81 40.98 ;
      RECT 160.47 38.7 160.63 40.98 ;
      RECT 160.47 40.03 160.81 40.31 ;
      RECT 160.47 38.7 160.81 38.98 ;
      RECT 160.11 55.68 160.27 56.51 ;
      RECT 159.87 55.68 160.27 55.84 ;
      RECT 159.87 53.67 160.03 55.84 ;
      RECT 159.87 53.67 160.51 53.83 ;
      RECT 160.23 53.35 160.51 53.83 ;
      RECT 159.97 51.7 160.35 51.92 ;
      RECT 160.19 50.98 160.35 51.92 ;
      RECT 159.55 52.58 160.31 52.86 ;
      RECT 160.15 52.18 160.31 52.86 ;
      RECT 159.55 51.64 159.71 52.86 ;
      RECT 159.87 62.9 160.03 67.89 ;
      RECT 159.87 65.82 160.09 66.55 ;
      RECT 159.55 47.39 159.71 49.72 ;
      RECT 159.55 47.39 160.03 47.55 ;
      RECT 159.87 43.85 160.03 47.55 ;
      RECT 159.25 43.85 160.03 44.01 ;
      RECT 159.25 39.56 159.41 44.01 ;
      RECT 159.25 39.56 159.59 39.84 ;
      RECT 159.43 39.16 159.59 39.84 ;
      RECT 159.57 34.44 159.91 34.72 ;
      RECT 159.75 32.44 159.91 34.72 ;
      RECT 159.57 33.11 159.91 33.39 ;
      RECT 159.57 32.44 159.91 32.72 ;
      RECT 159.57 40.7 159.91 40.98 ;
      RECT 159.75 38.7 159.91 40.98 ;
      RECT 159.57 40.03 159.91 40.31 ;
      RECT 159.57 38.7 159.91 38.98 ;
      RECT 159.39 62.9 159.55 67.89 ;
      RECT 159.39 64.59 159.67 65.31 ;
      RECT 158.91 46.75 159.07 47.43 ;
      RECT 158.59 46.75 159.39 46.91 ;
      RECT 159.23 44.23 159.39 46.91 ;
      RECT 158.59 44.23 158.75 46.91 ;
      RECT 156.69 34.88 158.89 35.04 ;
      RECT 158.61 34.59 158.89 35.04 ;
      RECT 157.67 34.59 157.91 35.04 ;
      RECT 156.69 34.59 156.97 35.04 ;
      RECT 157.67 38.38 157.91 39.02 ;
      RECT 158.61 38.38 158.89 38.83 ;
      RECT 156.69 38.38 156.97 38.83 ;
      RECT 156.69 38.38 158.89 38.54 ;
      RECT 156.85 36.47 158.73 36.63 ;
      RECT 158.57 35.88 158.73 36.63 ;
      RECT 157.71 35.23 157.87 36.63 ;
      RECT 156.85 35.88 157.01 36.63 ;
      RECT 158.67 35.23 158.83 36.06 ;
      RECT 156.75 35.23 156.91 36.06 ;
      RECT 158.67 37.11 158.83 38.19 ;
      RECT 157.71 36.79 157.87 38.19 ;
      RECT 156.75 37.11 156.91 38.19 ;
      RECT 158.57 36.79 158.73 37.39 ;
      RECT 156.85 36.79 157.01 37.39 ;
      RECT 156.85 36.79 158.73 36.95 ;
      RECT 156.93 68.07 158.75 68.23 ;
      RECT 156.93 62.02 157.09 68.23 ;
      RECT 156.93 62.02 157.31 62.18 ;
      RECT 157.15 57.45 157.31 62.18 ;
      RECT 157.15 57.45 158.75 57.61 ;
      RECT 158.43 57.39 158.75 57.61 ;
      RECT 158.43 53.74 158.59 57.61 ;
      RECT 158.59 51.32 158.75 53.9 ;
      RECT 158.27 51.32 158.75 51.48 ;
      RECT 158.27 49.88 158.43 51.48 ;
      RECT 157.95 49.88 158.43 50.04 ;
      RECT 157.95 47.71 158.11 50.04 ;
      RECT 157.49 47.71 158.11 47.99 ;
      RECT 158.27 47.39 158.43 49.72 ;
      RECT 157.95 47.39 158.43 47.55 ;
      RECT 157.95 43.85 158.11 47.55 ;
      RECT 157.95 43.85 158.73 44.01 ;
      RECT 158.57 39.56 158.73 44.01 ;
      RECT 158.39 39.56 158.73 39.84 ;
      RECT 158.39 39.16 158.55 39.84 ;
      RECT 158.43 62.9 158.59 67.89 ;
      RECT 158.31 64.59 158.59 65.31 ;
      RECT 157.67 52.58 158.43 52.86 ;
      RECT 158.27 51.64 158.43 52.86 ;
      RECT 157.67 52.18 157.83 52.86 ;
      RECT 158.07 34.44 158.41 34.72 ;
      RECT 158.07 32.44 158.23 34.72 ;
      RECT 158.07 33.11 158.41 33.39 ;
      RECT 158.07 32.44 158.41 32.72 ;
      RECT 158.07 40.7 158.41 40.98 ;
      RECT 158.07 38.7 158.23 40.98 ;
      RECT 158.07 40.03 158.41 40.31 ;
      RECT 158.07 38.7 158.41 38.98 ;
      RECT 158.13 53.23 158.41 53.51 ;
      RECT 158.13 53.03 158.29 53.51 ;
      RECT 157.31 53.03 158.29 53.19 ;
      RECT 157.31 50.98 157.47 53.19 ;
      RECT 157.27 52.54 157.47 52.82 ;
      RECT 156.93 50.98 157.47 51.14 ;
      RECT 156.93 50.8 157.15 51.14 ;
      RECT 156.83 56.67 156.99 61.86 ;
      RECT 156.83 56.67 158.27 56.83 ;
      RECT 158.11 56 158.27 56.83 ;
      RECT 156.99 54.4 157.15 56.83 ;
      RECT 157.95 50.66 158.11 51.5 ;
      RECT 157.31 50.66 158.11 50.82 ;
      RECT 157.31 50.18 157.47 50.82 ;
      RECT 156.83 50.18 157.47 50.5 ;
      RECT 156.83 47.07 156.99 50.5 ;
      RECT 156.83 47.07 157.31 47.23 ;
      RECT 157.15 45.44 157.31 47.23 ;
      RECT 157.71 55.68 157.87 56.51 ;
      RECT 157.71 55.68 158.11 55.84 ;
      RECT 157.95 53.67 158.11 55.84 ;
      RECT 157.47 53.67 158.11 53.83 ;
      RECT 157.47 53.35 157.75 53.83 ;
      RECT 157.95 62.9 158.11 67.89 ;
      RECT 157.89 65.82 158.11 66.55 ;
      RECT 157.63 51.7 158.01 51.92 ;
      RECT 157.63 50.98 157.79 51.92 ;
      RECT 157.15 47.39 157.31 49.72 ;
      RECT 157.15 47.39 157.63 47.55 ;
      RECT 157.47 43.85 157.63 47.55 ;
      RECT 156.85 43.85 157.63 44.01 ;
      RECT 156.85 39.56 157.01 44.01 ;
      RECT 156.85 39.56 157.19 39.84 ;
      RECT 157.03 39.16 157.19 39.84 ;
      RECT 157.17 34.44 157.51 34.72 ;
      RECT 157.35 32.44 157.51 34.72 ;
      RECT 157.17 33.11 157.51 33.39 ;
      RECT 157.17 32.44 157.51 32.72 ;
      RECT 157.17 40.7 157.51 40.98 ;
      RECT 157.35 38.7 157.51 40.98 ;
      RECT 157.17 40.03 157.51 40.31 ;
      RECT 157.17 38.7 157.51 38.98 ;
      RECT 157.31 54.06 157.47 56.51 ;
      RECT 156.95 54.06 157.47 54.22 ;
      RECT 156.95 52.98 157.15 54.22 ;
      RECT 156.95 51.34 157.11 54.22 ;
      RECT 156.95 51.34 157.15 52.12 ;
      RECT 156.51 46.75 156.67 47.43 ;
      RECT 156.19 46.75 156.99 46.91 ;
      RECT 156.83 44.23 156.99 46.91 ;
      RECT 156.19 44.23 156.35 46.91 ;
      RECT 154.29 34.88 156.49 35.04 ;
      RECT 156.21 34.59 156.49 35.04 ;
      RECT 155.27 34.59 155.51 35.04 ;
      RECT 154.29 34.59 154.57 35.04 ;
      RECT 155.27 38.38 155.51 39.02 ;
      RECT 156.21 38.38 156.49 38.83 ;
      RECT 154.29 38.38 154.57 38.83 ;
      RECT 154.29 38.38 156.49 38.54 ;
      RECT 154.45 36.47 156.33 36.63 ;
      RECT 156.17 35.86 156.33 36.63 ;
      RECT 155.31 35.23 155.47 36.63 ;
      RECT 154.45 35.86 154.61 36.63 ;
      RECT 156.27 35.23 156.43 36.05 ;
      RECT 154.35 35.23 154.51 36.05 ;
      RECT 156.27 37.11 156.43 38.19 ;
      RECT 155.31 36.79 155.47 38.19 ;
      RECT 154.35 37.11 154.51 38.19 ;
      RECT 156.17 36.79 156.33 37.39 ;
      RECT 154.45 36.79 154.61 37.39 ;
      RECT 154.45 36.79 156.33 36.95 ;
      RECT 155.07 50.66 155.23 51.5 ;
      RECT 155.07 50.66 155.87 50.82 ;
      RECT 155.71 50.18 155.87 50.82 ;
      RECT 155.71 50.18 156.35 50.5 ;
      RECT 156.19 47.07 156.35 50.5 ;
      RECT 155.87 47.07 156.35 47.23 ;
      RECT 155.87 45.44 156.03 47.23 ;
      RECT 156.19 56.67 156.35 61.86 ;
      RECT 154.91 56.67 156.35 56.83 ;
      RECT 156.03 54.4 156.19 56.83 ;
      RECT 154.91 56 155.07 56.83 ;
      RECT 155.87 47.39 156.03 49.72 ;
      RECT 155.55 47.39 156.03 47.55 ;
      RECT 155.55 43.85 155.71 47.55 ;
      RECT 155.55 43.85 156.33 44.01 ;
      RECT 156.17 39.56 156.33 44.01 ;
      RECT 155.99 39.56 156.33 39.84 ;
      RECT 155.99 39.16 156.15 39.84 ;
      RECT 154.77 53.23 155.05 53.51 ;
      RECT 154.89 53.03 155.05 53.51 ;
      RECT 154.89 53.03 155.87 53.19 ;
      RECT 155.71 50.98 155.87 53.19 ;
      RECT 155.71 52.54 155.91 52.82 ;
      RECT 155.71 50.98 156.25 51.14 ;
      RECT 156.03 50.8 156.25 51.14 ;
      RECT 154.43 68.07 156.25 68.23 ;
      RECT 156.09 62.02 156.25 68.23 ;
      RECT 155.87 62.02 156.25 62.18 ;
      RECT 155.87 57.45 156.03 62.18 ;
      RECT 154.43 57.45 156.03 57.61 ;
      RECT 154.43 57.39 154.75 57.61 ;
      RECT 154.59 53.74 154.75 57.61 ;
      RECT 154.43 51.32 154.59 53.9 ;
      RECT 154.43 51.32 154.91 51.48 ;
      RECT 154.75 49.88 154.91 51.48 ;
      RECT 154.75 49.88 155.23 50.04 ;
      RECT 155.07 47.71 155.23 50.04 ;
      RECT 155.07 47.71 155.69 47.99 ;
      RECT 155.71 54.06 155.87 56.51 ;
      RECT 155.71 54.06 156.23 54.22 ;
      RECT 156.07 51.34 156.23 54.22 ;
      RECT 156.03 52.98 156.23 54.22 ;
      RECT 156.03 51.34 156.23 52.12 ;
      RECT 155.67 34.44 156.01 34.72 ;
      RECT 155.67 32.44 155.83 34.72 ;
      RECT 155.67 33.11 156.01 33.39 ;
      RECT 155.67 32.44 156.01 32.72 ;
      RECT 155.67 40.7 156.01 40.98 ;
      RECT 155.67 38.7 155.83 40.98 ;
      RECT 155.67 40.03 156.01 40.31 ;
      RECT 155.67 38.7 156.01 38.98 ;
      RECT 155.31 55.68 155.47 56.51 ;
      RECT 155.07 55.68 155.47 55.84 ;
      RECT 155.07 53.67 155.23 55.84 ;
      RECT 155.07 53.67 155.71 53.83 ;
      RECT 155.43 53.35 155.71 53.83 ;
      RECT 155.17 51.7 155.55 51.92 ;
      RECT 155.39 50.98 155.55 51.92 ;
      RECT 154.75 52.58 155.51 52.86 ;
      RECT 155.35 52.18 155.51 52.86 ;
      RECT 154.75 51.64 154.91 52.86 ;
      RECT 155.07 62.9 155.23 67.89 ;
      RECT 155.07 65.82 155.29 66.55 ;
      RECT 154.75 47.39 154.91 49.72 ;
      RECT 154.75 47.39 155.23 47.55 ;
      RECT 155.07 43.85 155.23 47.55 ;
      RECT 154.45 43.85 155.23 44.01 ;
      RECT 154.45 39.56 154.61 44.01 ;
      RECT 154.45 39.56 154.79 39.84 ;
      RECT 154.63 39.16 154.79 39.84 ;
      RECT 154.77 34.44 155.11 34.72 ;
      RECT 154.95 32.44 155.11 34.72 ;
      RECT 154.77 33.11 155.11 33.39 ;
      RECT 154.77 32.44 155.11 32.72 ;
      RECT 154.77 40.7 155.11 40.98 ;
      RECT 154.95 38.7 155.11 40.98 ;
      RECT 154.77 40.03 155.11 40.31 ;
      RECT 154.77 38.7 155.11 38.98 ;
      RECT 154.59 62.9 154.75 67.89 ;
      RECT 154.59 64.59 154.87 65.31 ;
      RECT 154.11 46.75 154.27 47.43 ;
      RECT 154.11 46.75 154.59 46.91 ;
      RECT 154.43 44.23 154.59 46.91 ;
      RECT 149.74 12.78 153.62 14.94 ;
      RECT 142.31 13.62 153.62 14.18 ;
      RECT 142.31 10.25 142.87 14.18 ;
      RECT 151.04 10.15 152.58 14.94 ;
      RECT 142.31 11.93 146.2 12.49 ;
      RECT 149.05 11.46 149.33 11.62 ;
      RECT 151.04 10.15 153.32 11.51 ;
      RECT 149.11 10.25 149.27 11.62 ;
      RECT 141.5 10.25 149.27 10.81 ;
      RECT 152.13 30.09 152.29 43.81 ;
      RECT 152.13 30.09 153.39 30.25 ;
      RECT 153.23 16.21 153.39 30.25 ;
      RECT 150.69 68.06 153.29 68.66 ;
      RECT 153.09 67.94 153.29 68.66 ;
      RECT 151.29 39.38 151.45 68.66 ;
      RECT 152.91 16.98 153.07 24 ;
      RECT 151.85 16.98 153.07 17.14 ;
      RECT 151.45 29.77 153.03 29.93 ;
      RECT 152.87 29.42 153.03 29.93 ;
      RECT 152.41 26.46 152.57 29.93 ;
      RECT 151.45 26.46 151.61 29.93 ;
      RECT 150.99 28.06 151.61 29.16 ;
      RECT 151.93 25.88 152.09 29.61 ;
      RECT 151.93 25.88 152.75 26.04 ;
      RECT 152.59 21.53 152.75 26.04 ;
      RECT 151.21 21.53 152.75 21.69 ;
      RECT 151.21 21.16 151.37 21.69 ;
      RECT 150.09 21.16 151.37 21.32 ;
      RECT 151.05 18.36 151.21 21.32 ;
      RECT 150.09 18.36 150.25 21.32 ;
      RECT 143.57 25.85 151.35 26.01 ;
      RECT 151.19 25.56 151.35 26.01 ;
      RECT 151.19 25.56 152.43 25.72 ;
      RECT 152.27 22.17 152.43 25.72 ;
      RECT 150.31 22.81 151.21 22.97 ;
      RECT 151.05 22.17 151.21 22.97 ;
      RECT 150.31 21.97 150.47 22.97 ;
      RECT 151.05 22.17 152.43 22.33 ;
      RECT 148.33 21.97 150.47 22.13 ;
      RECT 149.13 18.36 149.29 22.13 ;
      RECT 148.33 21.45 148.49 22.13 ;
      RECT 151.53 17.29 151.69 21.37 ;
      RECT 149.61 17.49 149.77 21.19 ;
      RECT 150.57 17.73 150.73 21 ;
      RECT 152.17 17.73 152.33 18.26 ;
      RECT 149.61 17.73 152.33 17.91 ;
      RECT 151.49 17.29 151.69 17.91 ;
      RECT 150.41 17.29 150.57 17.91 ;
      RECT 151.35 30.63 151.55 32.75 ;
      RECT 151.35 31.81 151.97 32.09 ;
      RECT 150.89 35.36 151.21 35.52 ;
      RECT 151.05 32.97 151.21 35.52 ;
      RECT 151.05 32.97 151.89 33.13 ;
      RECT 151.73 32.38 151.89 33.13 ;
      RECT 150.85 30.29 151.53 30.45 ;
      RECT 150.85 29.48 151.01 30.45 ;
      RECT 150.85 29.48 151.17 29.64 ;
      RECT 150.87 30.63 151.03 32.75 ;
      RECT 150.53 30.63 151.03 30.79 ;
      RECT 150.53 26.85 150.69 30.79 ;
      RECT 150.53 26.85 151.21 27.01 ;
      RECT 151.05 26.19 151.21 27.01 ;
      RECT 150.97 16.95 151.13 17.57 ;
      RECT 150.61 16.95 151.13 17.11 ;
      RECT 150.61 15.3 150.77 17.11 ;
      RECT 148.59 15.3 150.77 15.46 ;
      RECT 143.83 25.53 151.03 25.69 ;
      RECT 150.87 23.88 151.03 25.69 ;
      RECT 149.11 23.88 149.27 25.69 ;
      RECT 147.35 22.06 147.51 25.69 ;
      RECT 145.59 17.87 145.75 25.69 ;
      RECT 143.83 23.78 143.99 25.69 ;
      RECT 145.59 22.06 148.13 22.22 ;
      RECT 147.97 18.97 148.13 22.22 ;
      RECT 146.55 17.87 146.71 22.22 ;
      RECT 150.73 21.48 150.89 22.65 ;
      RECT 149.83 21.48 150.91 21.69 ;
      RECT 150.51 33.79 150.67 36.17 ;
      RECT 148.59 33.79 148.75 36.17 ;
      RECT 146.67 33.79 146.83 36.17 ;
      RECT 144.75 33.79 144.91 36.17 ;
      RECT 142.83 33.79 142.99 36.17 ;
      RECT 140.91 33.79 141.07 36.17 ;
      RECT 149.55 34.1 149.71 34.66 ;
      RECT 147.63 34.1 147.79 34.66 ;
      RECT 145.71 34.1 145.87 34.66 ;
      RECT 143.79 34.1 143.95 34.66 ;
      RECT 141.87 34.1 142.03 34.66 ;
      RECT 140.91 34.1 150.67 34.26 ;
      RECT 150.51 36.4 150.67 42.37 ;
      RECT 149.55 37.67 149.71 42.37 ;
      RECT 148.59 36.4 148.75 42.37 ;
      RECT 147.63 37.67 147.79 42.37 ;
      RECT 146.67 36.4 146.83 42.37 ;
      RECT 145.71 37.67 145.87 42.37 ;
      RECT 144.75 36.4 144.91 42.37 ;
      RECT 143.79 37.67 143.95 42.37 ;
      RECT 142.83 36.4 142.99 42.37 ;
      RECT 141.87 37.67 142.03 42.37 ;
      RECT 140.91 36.4 141.07 42.37 ;
      RECT 140.91 37.67 150.67 37.83 ;
      RECT 149.55 36.87 150.67 37.03 ;
      RECT 145.71 36.87 147.79 37.03 ;
      RECT 147.63 36.4 147.79 37.03 ;
      RECT 141.87 36.87 143.95 37.03 ;
      RECT 143.79 36.4 143.95 37.03 ;
      RECT 149.55 36.4 149.71 37.03 ;
      RECT 145.71 36.4 145.87 37.03 ;
      RECT 141.87 36.4 142.03 37.03 ;
      RECT 149.55 47.16 149.71 51.33 ;
      RECT 149.55 48.4 150.67 48.59 ;
      RECT 150.51 47.14 150.67 48.59 ;
      RECT 149.87 42.85 150.17 43.09 ;
      RECT 149.87 42.85 150.45 43.03 ;
      RECT 148.91 52.33 150.35 52.55 ;
      RECT 150.13 51.48 150.35 52.55 ;
      RECT 146.99 52.33 148.43 52.55 ;
      RECT 148.21 51.44 148.43 52.55 ;
      RECT 148.91 51.44 149.13 52.55 ;
      RECT 146.99 51.48 147.21 52.55 ;
      RECT 150.03 48.78 150.19 51.77 ;
      RECT 149.07 46.79 149.23 51.77 ;
      RECT 148.11 46.79 148.27 51.77 ;
      RECT 147.15 48.78 147.31 51.77 ;
      RECT 149.07 46.79 149.87 47 ;
      RECT 147.47 46.79 148.27 47 ;
      RECT 147.47 46.79 149.87 46.96 ;
      RECT 148.59 43.19 148.75 46.96 ;
      RECT 149.07 37.35 150.15 37.51 ;
      RECT 149.07 35.68 149.23 37.51 ;
      RECT 150.03 35.68 150.19 36.68 ;
      RECT 148.97 35.68 150.29 35.84 ;
      RECT 150.13 34.58 150.29 35.84 ;
      RECT 148.97 34.58 149.13 35.84 ;
      RECT 150.03 34.58 150.29 34.86 ;
      RECT 148.97 34.58 149.23 34.86 ;
      RECT 149.55 42.53 149.71 46.23 ;
      RECT 149.07 42.53 150.19 42.69 ;
      RECT 150.03 37.99 150.19 42.69 ;
      RECT 149.07 37.99 149.23 42.69 ;
      RECT 150.03 43.34 150.19 47.95 ;
      RECT 149.07 46.47 150.19 46.63 ;
      RECT 149.07 43.34 149.23 46.63 ;
      RECT 148.77 18.02 149.45 18.18 ;
      RECT 149.29 16.98 149.45 18.18 ;
      RECT 149.29 16.98 150.15 17.14 ;
      RECT 148.91 33.1 150.03 33.26 ;
      RECT 149.87 30.63 150.03 33.26 ;
      RECT 148.91 30.63 149.07 33.26 ;
      RECT 149.29 51.95 149.97 52.11 ;
      RECT 149.55 51.6 149.71 52.11 ;
      RECT 146.09 510.04 147.41 510.94 ;
      RECT 142.25 510.04 143.57 510.94 ;
      RECT 135.01 510.04 137.81 510.94 ;
      RECT 128.21 510.04 131.01 510.94 ;
      RECT 121.41 510.04 124.21 510.94 ;
      RECT 114.61 510.04 117.41 510.94 ;
      RECT 109.51 510.04 110.61 510.94 ;
      RECT 106.11 510.04 107.21 510.94 ;
      RECT 102.71 510.04 103.81 510.94 ;
      RECT 99.31 510.04 100.41 510.94 ;
      RECT 95.91 510.04 97.01 510.94 ;
      RECT 92.51 510.04 93.61 510.94 ;
      RECT 89.11 510.04 90.21 510.94 ;
      RECT 86.61 510.04 87.41 510.94 ;
      RECT 85.41 510.04 86.21 510.94 ;
      RECT 81.81 510.04 82.61 510.94 ;
      RECT 80.61 510.04 81.41 510.94 ;
      RECT 77.01 510.04 77.81 510.94 ;
      RECT 75.81 510.04 76.61 510.94 ;
      RECT 72.21 510.04 73.01 510.94 ;
      RECT 71.01 510.04 71.81 510.94 ;
      RECT 67.41 510.04 68.21 510.94 ;
      RECT 66.21 510.04 67.01 510.94 ;
      RECT 62.61 510.04 63.41 510.94 ;
      RECT 61.41 510.04 62.21 510.94 ;
      RECT 57.81 510.04 58.61 510.94 ;
      RECT 56.61 510.04 57.41 510.94 ;
      RECT 53.01 510.04 53.81 510.94 ;
      RECT 51.81 510.04 52.61 510.94 ;
      RECT 48.21 510.04 49.01 510.94 ;
      RECT 47.01 510.04 47.81 510.94 ;
      RECT 45.81 510.04 46.61 510.94 ;
      RECT 42.21 510.04 43.01 510.94 ;
      RECT 41.01 510.04 41.81 510.94 ;
      RECT 37.41 510.04 38.21 510.94 ;
      RECT 36.21 510.04 37.01 510.94 ;
      RECT 32.61 510.04 33.41 510.94 ;
      RECT 31.41 510.04 32.21 510.94 ;
      RECT 27.81 510.04 28.61 510.94 ;
      RECT 26.61 510.04 27.41 510.94 ;
      RECT 23.01 510.04 23.81 510.94 ;
      RECT 21.81 510.04 22.61 510.94 ;
      RECT 18.21 510.04 19.01 510.94 ;
      RECT 17.01 510.04 17.81 510.94 ;
      RECT 13.41 510.04 14.21 510.94 ;
      RECT 12.21 510.04 13.01 510.94 ;
      RECT 8.61 510.04 9.41 510.94 ;
      RECT 7.41 510.04 8.21 510.94 ;
      RECT 85.41 510.04 87.41 510.74 ;
      RECT 80.61 510.04 82.61 510.74 ;
      RECT 75.81 510.04 77.81 510.74 ;
      RECT 71.01 510.04 73.01 510.74 ;
      RECT 66.21 510.04 68.21 510.74 ;
      RECT 61.41 510.04 63.41 510.74 ;
      RECT 56.61 510.04 58.61 510.74 ;
      RECT 51.81 510.04 53.81 510.74 ;
      RECT 45.81 510.04 49.01 510.74 ;
      RECT 41.01 510.04 43.01 510.74 ;
      RECT 36.21 510.04 38.21 510.74 ;
      RECT 31.41 510.04 33.41 510.74 ;
      RECT 26.61 510.04 28.61 510.74 ;
      RECT 21.81 510.04 23.81 510.74 ;
      RECT 17.01 510.04 19.01 510.74 ;
      RECT 12.21 510.04 14.21 510.74 ;
      RECT 7.21 510.04 9.41 510.74 ;
      RECT 7.21 510.04 87.41 510.22 ;
      RECT 6.98 510.04 149.93 510.2 ;
      RECT 149.77 69.48 149.93 510.2 ;
      RECT 85.73 68.88 85.89 510.94 ;
      RECT 84.53 68.88 84.69 510.22 ;
      RECT 83.33 68.88 83.49 510.22 ;
      RECT 82.13 68.88 82.29 510.94 ;
      RECT 80.93 68.88 81.09 510.94 ;
      RECT 79.73 68.88 79.89 510.22 ;
      RECT 78.53 68.88 78.69 510.22 ;
      RECT 77.33 68.88 77.49 510.94 ;
      RECT 76.13 68.88 76.29 510.94 ;
      RECT 74.93 68.88 75.09 510.22 ;
      RECT 73.73 68.88 73.89 510.22 ;
      RECT 72.53 68.88 72.69 510.94 ;
      RECT 71.33 68.88 71.49 510.94 ;
      RECT 70.13 68.88 70.29 510.22 ;
      RECT 68.93 68.88 69.09 510.22 ;
      RECT 67.73 68.88 67.89 510.94 ;
      RECT 66.53 68.88 66.69 510.94 ;
      RECT 65.33 68.88 65.49 510.22 ;
      RECT 64.13 68.88 64.29 510.22 ;
      RECT 62.93 68.88 63.09 510.94 ;
      RECT 61.73 68.88 61.89 510.94 ;
      RECT 60.53 68.88 60.69 510.22 ;
      RECT 59.33 68.88 59.49 510.22 ;
      RECT 58.13 68.88 58.29 510.94 ;
      RECT 56.93 68.88 57.09 510.94 ;
      RECT 55.73 68.88 55.89 510.22 ;
      RECT 54.53 68.88 54.69 510.22 ;
      RECT 53.33 68.88 53.49 510.94 ;
      RECT 52.13 68.88 52.29 510.94 ;
      RECT 50.93 68.88 51.09 510.22 ;
      RECT 49.73 68.88 49.89 510.22 ;
      RECT 48.53 68.88 48.69 510.94 ;
      RECT 46.13 68.88 46.29 510.94 ;
      RECT 44.93 68.88 45.09 510.22 ;
      RECT 43.73 68.88 43.89 510.22 ;
      RECT 42.53 68.88 42.69 510.94 ;
      RECT 41.33 68.88 41.49 510.94 ;
      RECT 40.13 68.88 40.29 510.22 ;
      RECT 38.93 68.88 39.09 510.22 ;
      RECT 37.73 68.88 37.89 510.94 ;
      RECT 36.53 68.88 36.69 510.94 ;
      RECT 35.33 68.88 35.49 510.22 ;
      RECT 34.13 68.88 34.29 510.22 ;
      RECT 32.93 68.88 33.09 510.94 ;
      RECT 31.73 68.88 31.89 510.94 ;
      RECT 30.53 68.88 30.69 510.22 ;
      RECT 29.33 68.88 29.49 510.22 ;
      RECT 28.13 68.88 28.29 510.94 ;
      RECT 26.93 68.88 27.09 510.94 ;
      RECT 25.73 68.88 25.89 510.22 ;
      RECT 24.53 68.88 24.69 510.22 ;
      RECT 23.33 68.88 23.49 510.94 ;
      RECT 22.13 68.88 22.29 510.94 ;
      RECT 20.93 68.88 21.09 510.22 ;
      RECT 19.73 68.88 19.89 510.22 ;
      RECT 18.53 68.88 18.69 510.94 ;
      RECT 17.33 68.88 17.49 510.94 ;
      RECT 16.13 68.88 16.29 510.22 ;
      RECT 14.93 68.88 15.09 510.22 ;
      RECT 13.73 68.88 13.89 510.94 ;
      RECT 12.53 68.88 12.69 510.94 ;
      RECT 11.33 68.88 11.49 510.22 ;
      RECT 10.13 68.88 10.29 510.22 ;
      RECT 8.93 68.88 9.09 510.94 ;
      RECT 6.98 67.81 7.14 510.2 ;
      RECT 7.38 68.88 87.44 509.88 ;
      RECT 6.98 509.46 87.68 509.69 ;
      RECT 7.38 509.03 88.22 509.3 ;
      RECT 87.71 505.7 87.89 509.3 ;
      RECT 6.24 506.6 7.14 508.6 ;
      RECT 7.38 505.7 88.22 505.97 ;
      RECT 145.22 505.64 149.93 505.8 ;
      RECT 6.98 505.2 87.61 505.36 ;
      RECT 7.38 504.59 88.22 504.86 ;
      RECT 144.63 504.68 149.93 504.84 ;
      RECT 87.71 69.46 87.89 504.86 ;
      RECT 145.22 503.72 149.93 503.88 ;
      RECT 6.24 502.66 7.14 503.46 ;
      RECT 149.63 502.72 149.93 503.42 ;
      RECT 145.22 502.24 149.93 502.4 ;
      RECT 7.38 501.19 88.22 501.53 ;
      RECT 144.57 501.28 149.93 501.44 ;
      RECT 145.22 500.32 149.93 500.48 ;
      RECT 6.24 499.26 7.14 500.06 ;
      RECT 149.63 499.3 149.93 500 ;
      RECT 145.22 498.84 149.93 499 ;
      RECT 7.38 497.79 88.22 498.13 ;
      RECT 144.63 497.88 149.93 498.04 ;
      RECT 145.22 496.92 149.93 497.08 ;
      RECT 6.24 495.86 7.14 496.66 ;
      RECT 149.63 495.92 149.93 496.62 ;
      RECT 145.22 495.44 149.93 495.6 ;
      RECT 7.38 494.39 88.22 494.73 ;
      RECT 144.57 494.48 149.93 494.64 ;
      RECT 145.22 493.52 149.93 493.68 ;
      RECT 6.24 492.46 7.14 493.26 ;
      RECT 149.63 492.5 149.93 493.2 ;
      RECT 145.22 492.04 149.93 492.2 ;
      RECT 7.38 490.99 88.22 491.33 ;
      RECT 144.63 491.08 149.93 491.24 ;
      RECT 145.22 490.12 149.93 490.28 ;
      RECT 6.24 489.06 7.14 489.86 ;
      RECT 149.63 489.12 149.93 489.82 ;
      RECT 145.22 488.64 149.93 488.8 ;
      RECT 7.38 487.59 88.22 487.93 ;
      RECT 144.57 487.68 149.93 487.84 ;
      RECT 145.22 486.72 149.93 486.88 ;
      RECT 6.24 485.66 7.14 486.46 ;
      RECT 149.63 485.7 149.93 486.4 ;
      RECT 145.22 485.24 149.93 485.4 ;
      RECT 7.38 484.19 88.22 484.53 ;
      RECT 144.63 484.28 149.93 484.44 ;
      RECT 145.22 483.32 149.93 483.48 ;
      RECT 6.24 482.26 7.14 483.06 ;
      RECT 149.63 482.32 149.93 483.02 ;
      RECT 145.22 481.84 149.93 482 ;
      RECT 7.38 480.79 88.22 481.13 ;
      RECT 144.57 480.88 149.93 481.04 ;
      RECT 145.22 479.92 149.93 480.08 ;
      RECT 6.24 478.86 7.14 479.66 ;
      RECT 149.63 478.9 149.93 479.6 ;
      RECT 145.22 478.44 149.93 478.6 ;
      RECT 7.38 477.39 88.22 477.73 ;
      RECT 144.63 477.48 149.93 477.64 ;
      RECT 145.22 476.52 149.93 476.68 ;
      RECT 6.24 475.46 7.14 476.26 ;
      RECT 149.63 475.52 149.93 476.22 ;
      RECT 145.22 475.04 149.93 475.2 ;
      RECT 7.38 473.99 88.22 474.33 ;
      RECT 144.57 474.08 149.93 474.24 ;
      RECT 145.22 473.12 149.93 473.28 ;
      RECT 6.24 472.06 7.14 472.86 ;
      RECT 149.63 472.1 149.93 472.8 ;
      RECT 145.22 471.64 149.93 471.8 ;
      RECT 7.38 470.59 88.22 470.93 ;
      RECT 144.63 470.68 149.93 470.84 ;
      RECT 145.22 469.72 149.93 469.88 ;
      RECT 6.24 468.66 7.14 469.46 ;
      RECT 149.63 468.72 149.93 469.42 ;
      RECT 145.22 468.24 149.93 468.4 ;
      RECT 7.38 467.19 88.22 467.53 ;
      RECT 144.57 467.28 149.93 467.44 ;
      RECT 145.22 466.32 149.93 466.48 ;
      RECT 6.24 465.26 7.14 466.06 ;
      RECT 149.63 465.3 149.93 466 ;
      RECT 145.22 464.84 149.93 465 ;
      RECT 7.38 463.79 88.22 464.13 ;
      RECT 144.63 463.88 149.93 464.04 ;
      RECT 145.22 462.92 149.93 463.08 ;
      RECT 6.24 461.86 7.14 462.66 ;
      RECT 149.63 461.92 149.93 462.62 ;
      RECT 145.22 461.44 149.93 461.6 ;
      RECT 7.38 460.39 88.22 460.73 ;
      RECT 144.57 460.48 149.93 460.64 ;
      RECT 145.22 459.52 149.93 459.68 ;
      RECT 6.24 458.46 7.14 459.26 ;
      RECT 149.63 458.5 149.93 459.2 ;
      RECT 145.22 458.04 149.93 458.2 ;
      RECT 7.38 456.99 88.22 457.33 ;
      RECT 144.63 457.08 149.93 457.24 ;
      RECT 145.22 456.12 149.93 456.28 ;
      RECT 6.24 455.06 7.14 455.86 ;
      RECT 149.63 455.12 149.93 455.82 ;
      RECT 145.22 454.64 149.93 454.8 ;
      RECT 7.38 453.59 88.22 453.93 ;
      RECT 144.57 453.68 149.93 453.84 ;
      RECT 145.22 452.72 149.93 452.88 ;
      RECT 6.24 451.66 7.14 452.46 ;
      RECT 149.63 451.7 149.93 452.4 ;
      RECT 145.22 451.24 149.93 451.4 ;
      RECT 7.38 450.19 88.22 450.53 ;
      RECT 144.63 450.28 149.93 450.44 ;
      RECT 145.22 449.32 149.93 449.48 ;
      RECT 6.24 448.26 7.14 449.06 ;
      RECT 149.63 448.32 149.93 449.02 ;
      RECT 145.22 447.84 149.93 448 ;
      RECT 7.38 446.79 88.22 447.13 ;
      RECT 144.57 446.88 149.93 447.04 ;
      RECT 145.22 445.92 149.93 446.08 ;
      RECT 6.24 444.86 7.14 445.66 ;
      RECT 149.63 444.9 149.93 445.6 ;
      RECT 145.22 444.44 149.93 444.6 ;
      RECT 7.38 443.39 88.22 443.73 ;
      RECT 144.63 443.48 149.93 443.64 ;
      RECT 145.22 442.52 149.93 442.68 ;
      RECT 6.24 441.46 7.14 442.26 ;
      RECT 149.63 441.52 149.93 442.22 ;
      RECT 145.22 441.04 149.93 441.2 ;
      RECT 7.38 439.99 88.22 440.33 ;
      RECT 144.57 440.08 149.93 440.24 ;
      RECT 145.22 439.12 149.93 439.28 ;
      RECT 6.24 438.06 7.14 438.86 ;
      RECT 149.63 438.1 149.93 438.8 ;
      RECT 145.22 437.64 149.93 437.8 ;
      RECT 7.38 436.59 88.22 436.93 ;
      RECT 144.63 436.68 149.93 436.84 ;
      RECT 145.22 435.72 149.93 435.88 ;
      RECT 6.24 434.66 7.14 435.46 ;
      RECT 149.63 434.72 149.93 435.42 ;
      RECT 145.22 434.24 149.93 434.4 ;
      RECT 7.38 433.19 88.22 433.53 ;
      RECT 144.57 433.28 149.93 433.44 ;
      RECT 145.22 432.32 149.93 432.48 ;
      RECT 6.24 431.26 7.14 432.06 ;
      RECT 149.63 431.3 149.93 432 ;
      RECT 145.22 430.84 149.93 431 ;
      RECT 7.38 429.79 88.22 430.13 ;
      RECT 144.63 429.88 149.93 430.04 ;
      RECT 145.22 428.92 149.93 429.08 ;
      RECT 6.24 427.86 7.14 428.66 ;
      RECT 149.63 427.92 149.93 428.62 ;
      RECT 145.22 427.44 149.93 427.6 ;
      RECT 7.38 426.39 88.22 426.73 ;
      RECT 144.57 426.48 149.93 426.64 ;
      RECT 145.22 425.52 149.93 425.68 ;
      RECT 6.24 424.46 7.14 425.26 ;
      RECT 149.63 424.5 149.93 425.2 ;
      RECT 145.22 424.04 149.93 424.2 ;
      RECT 7.38 422.99 88.22 423.33 ;
      RECT 144.63 423.08 149.93 423.24 ;
      RECT 145.22 422.12 149.93 422.28 ;
      RECT 6.24 421.06 7.14 421.86 ;
      RECT 149.63 421.12 149.93 421.82 ;
      RECT 145.22 420.64 149.93 420.8 ;
      RECT 7.38 419.59 88.22 419.93 ;
      RECT 144.57 419.68 149.93 419.84 ;
      RECT 145.22 418.72 149.93 418.88 ;
      RECT 6.24 417.66 7.14 418.46 ;
      RECT 149.63 417.7 149.93 418.4 ;
      RECT 145.22 417.24 149.93 417.4 ;
      RECT 7.38 416.19 88.22 416.53 ;
      RECT 144.63 416.28 149.93 416.44 ;
      RECT 145.22 415.32 149.93 415.48 ;
      RECT 6.24 414.26 7.14 415.06 ;
      RECT 149.63 414.32 149.93 415.02 ;
      RECT 145.22 413.84 149.93 414 ;
      RECT 7.38 412.79 88.22 413.13 ;
      RECT 144.57 412.88 149.93 413.04 ;
      RECT 145.22 411.92 149.93 412.08 ;
      RECT 6.24 410.86 7.14 411.66 ;
      RECT 149.63 410.9 149.93 411.6 ;
      RECT 145.22 410.44 149.93 410.6 ;
      RECT 7.38 409.39 88.22 409.73 ;
      RECT 144.63 409.48 149.93 409.64 ;
      RECT 145.22 408.52 149.93 408.68 ;
      RECT 6.24 407.46 7.14 408.26 ;
      RECT 149.63 407.52 149.93 408.22 ;
      RECT 145.22 407.04 149.93 407.2 ;
      RECT 7.38 405.99 88.22 406.33 ;
      RECT 144.57 406.08 149.93 406.24 ;
      RECT 145.22 405.12 149.93 405.28 ;
      RECT 6.24 404.06 7.14 404.86 ;
      RECT 149.63 404.1 149.93 404.8 ;
      RECT 145.22 403.64 149.93 403.8 ;
      RECT 7.38 402.59 88.22 402.93 ;
      RECT 144.63 402.68 149.93 402.84 ;
      RECT 145.22 401.72 149.93 401.88 ;
      RECT 6.24 400.66 7.14 401.46 ;
      RECT 149.63 400.72 149.93 401.42 ;
      RECT 145.22 400.24 149.93 400.4 ;
      RECT 7.38 399.19 88.22 399.53 ;
      RECT 144.57 399.28 149.93 399.44 ;
      RECT 145.22 398.32 149.93 398.48 ;
      RECT 6.24 397.26 7.14 398.06 ;
      RECT 149.63 397.3 149.93 398 ;
      RECT 145.22 396.84 149.93 397 ;
      RECT 7.38 395.79 88.22 396.13 ;
      RECT 144.63 395.88 149.93 396.04 ;
      RECT 145.22 394.92 149.93 395.08 ;
      RECT 6.24 393.86 7.14 394.66 ;
      RECT 149.63 393.92 149.93 394.62 ;
      RECT 145.22 393.44 149.93 393.6 ;
      RECT 7.38 392.39 88.22 392.73 ;
      RECT 144.57 392.48 149.93 392.64 ;
      RECT 145.22 391.52 149.93 391.68 ;
      RECT 6.24 390.46 7.14 391.26 ;
      RECT 149.63 390.5 149.93 391.2 ;
      RECT 145.22 390.04 149.93 390.2 ;
      RECT 7.38 388.99 88.22 389.33 ;
      RECT 144.63 389.08 149.93 389.24 ;
      RECT 145.22 388.12 149.93 388.28 ;
      RECT 6.24 387.06 7.14 387.86 ;
      RECT 149.63 387.12 149.93 387.82 ;
      RECT 145.22 386.64 149.93 386.8 ;
      RECT 7.38 385.59 88.22 385.93 ;
      RECT 144.57 385.68 149.93 385.84 ;
      RECT 145.22 384.72 149.93 384.88 ;
      RECT 6.24 383.66 7.14 384.46 ;
      RECT 149.63 383.7 149.93 384.4 ;
      RECT 145.22 383.24 149.93 383.4 ;
      RECT 7.38 382.19 88.22 382.53 ;
      RECT 144.63 382.28 149.93 382.44 ;
      RECT 145.22 381.32 149.93 381.48 ;
      RECT 6.24 380.26 7.14 381.06 ;
      RECT 149.63 380.32 149.93 381.02 ;
      RECT 145.22 379.84 149.93 380 ;
      RECT 7.38 378.79 88.22 379.13 ;
      RECT 144.57 378.88 149.93 379.04 ;
      RECT 145.22 377.92 149.93 378.08 ;
      RECT 6.24 376.86 7.14 377.66 ;
      RECT 149.63 376.9 149.93 377.6 ;
      RECT 145.22 376.44 149.93 376.6 ;
      RECT 7.38 375.39 88.22 375.73 ;
      RECT 144.63 375.48 149.93 375.64 ;
      RECT 145.22 374.52 149.93 374.68 ;
      RECT 6.24 373.46 7.14 374.26 ;
      RECT 149.63 373.52 149.93 374.22 ;
      RECT 145.22 373.04 149.93 373.2 ;
      RECT 7.38 371.99 88.22 372.33 ;
      RECT 144.57 372.08 149.93 372.24 ;
      RECT 145.22 371.12 149.93 371.28 ;
      RECT 6.24 370.06 7.14 370.86 ;
      RECT 149.63 370.1 149.93 370.8 ;
      RECT 145.22 369.64 149.93 369.8 ;
      RECT 7.38 368.59 88.22 368.93 ;
      RECT 144.63 368.68 149.93 368.84 ;
      RECT 145.22 367.72 149.93 367.88 ;
      RECT 6.24 366.66 7.14 367.46 ;
      RECT 149.63 366.72 149.93 367.42 ;
      RECT 145.22 366.24 149.93 366.4 ;
      RECT 7.38 365.19 88.22 365.53 ;
      RECT 144.57 365.28 149.93 365.44 ;
      RECT 145.22 364.32 149.93 364.48 ;
      RECT 6.24 363.26 7.14 364.06 ;
      RECT 149.63 363.3 149.93 364 ;
      RECT 145.22 362.84 149.93 363 ;
      RECT 7.38 361.79 88.22 362.13 ;
      RECT 144.63 361.88 149.93 362.04 ;
      RECT 145.22 360.92 149.93 361.08 ;
      RECT 6.24 359.86 7.14 360.66 ;
      RECT 149.63 359.92 149.93 360.62 ;
      RECT 145.22 359.44 149.93 359.6 ;
      RECT 7.38 358.39 88.22 358.73 ;
      RECT 144.57 358.48 149.93 358.64 ;
      RECT 145.22 357.52 149.93 357.68 ;
      RECT 6.24 356.46 7.14 357.26 ;
      RECT 149.63 356.5 149.93 357.2 ;
      RECT 145.22 356.04 149.93 356.2 ;
      RECT 7.38 354.99 88.22 355.33 ;
      RECT 144.63 355.08 149.93 355.24 ;
      RECT 145.22 354.12 149.93 354.28 ;
      RECT 6.24 353.06 7.14 353.86 ;
      RECT 149.63 353.12 149.93 353.82 ;
      RECT 145.22 352.64 149.93 352.8 ;
      RECT 7.38 351.59 88.22 351.93 ;
      RECT 144.57 351.68 149.93 351.84 ;
      RECT 145.22 350.72 149.93 350.88 ;
      RECT 6.24 349.66 7.14 350.46 ;
      RECT 149.63 349.7 149.93 350.4 ;
      RECT 145.22 349.24 149.93 349.4 ;
      RECT 7.38 348.19 88.22 348.53 ;
      RECT 144.63 348.28 149.93 348.44 ;
      RECT 145.22 347.32 149.93 347.48 ;
      RECT 6.24 346.26 7.14 347.06 ;
      RECT 149.63 346.32 149.93 347.02 ;
      RECT 145.22 345.84 149.93 346 ;
      RECT 7.38 344.79 88.22 345.13 ;
      RECT 144.57 344.88 149.93 345.04 ;
      RECT 145.22 343.92 149.93 344.08 ;
      RECT 6.24 342.86 7.14 343.66 ;
      RECT 149.63 342.9 149.93 343.6 ;
      RECT 145.22 342.44 149.93 342.6 ;
      RECT 7.38 341.39 88.22 341.73 ;
      RECT 144.63 341.48 149.93 341.64 ;
      RECT 145.22 340.52 149.93 340.68 ;
      RECT 6.24 339.46 7.14 340.26 ;
      RECT 149.63 339.52 149.93 340.22 ;
      RECT 145.22 339.04 149.93 339.2 ;
      RECT 7.38 337.99 88.22 338.33 ;
      RECT 144.57 338.08 149.93 338.24 ;
      RECT 145.22 337.12 149.93 337.28 ;
      RECT 6.24 336.06 7.14 336.86 ;
      RECT 149.63 336.1 149.93 336.8 ;
      RECT 145.22 335.64 149.93 335.8 ;
      RECT 7.38 334.59 88.22 334.93 ;
      RECT 144.63 334.68 149.93 334.84 ;
      RECT 145.22 333.72 149.93 333.88 ;
      RECT 6.24 332.66 7.14 333.46 ;
      RECT 149.63 332.72 149.93 333.42 ;
      RECT 145.22 332.24 149.93 332.4 ;
      RECT 7.38 331.19 88.22 331.53 ;
      RECT 144.57 331.28 149.93 331.44 ;
      RECT 145.22 330.32 149.93 330.48 ;
      RECT 6.24 329.26 7.14 330.06 ;
      RECT 149.63 329.3 149.93 330 ;
      RECT 145.22 328.84 149.93 329 ;
      RECT 7.38 327.79 88.22 328.13 ;
      RECT 144.63 327.88 149.93 328.04 ;
      RECT 145.22 326.92 149.93 327.08 ;
      RECT 6.24 325.86 7.14 326.66 ;
      RECT 149.63 325.92 149.93 326.62 ;
      RECT 145.22 325.44 149.93 325.6 ;
      RECT 7.38 324.39 88.22 324.73 ;
      RECT 144.57 324.48 149.93 324.64 ;
      RECT 145.22 323.52 149.93 323.68 ;
      RECT 6.24 322.46 7.14 323.26 ;
      RECT 149.63 322.5 149.93 323.2 ;
      RECT 145.22 322.04 149.93 322.2 ;
      RECT 7.38 320.99 88.22 321.33 ;
      RECT 144.63 321.08 149.93 321.24 ;
      RECT 145.22 320.12 149.93 320.28 ;
      RECT 6.24 319.06 7.14 319.86 ;
      RECT 149.63 319.12 149.93 319.82 ;
      RECT 145.22 318.64 149.93 318.8 ;
      RECT 7.38 317.59 88.22 317.93 ;
      RECT 144.57 317.68 149.93 317.84 ;
      RECT 145.22 316.72 149.93 316.88 ;
      RECT 6.24 315.66 7.14 316.46 ;
      RECT 149.63 315.7 149.93 316.4 ;
      RECT 145.22 315.24 149.93 315.4 ;
      RECT 7.38 314.19 88.22 314.53 ;
      RECT 144.63 314.28 149.93 314.44 ;
      RECT 145.22 313.32 149.93 313.48 ;
      RECT 6.24 312.26 7.14 313.06 ;
      RECT 149.63 312.32 149.93 313.02 ;
      RECT 145.22 311.84 149.93 312 ;
      RECT 7.38 310.79 88.22 311.13 ;
      RECT 144.57 310.88 149.93 311.04 ;
      RECT 145.22 309.92 149.93 310.08 ;
      RECT 6.24 308.86 7.14 309.66 ;
      RECT 149.63 308.9 149.93 309.6 ;
      RECT 145.22 308.44 149.93 308.6 ;
      RECT 7.38 307.39 88.22 307.73 ;
      RECT 144.63 307.48 149.93 307.64 ;
      RECT 145.22 306.52 149.93 306.68 ;
      RECT 6.24 305.46 7.14 306.26 ;
      RECT 149.63 305.52 149.93 306.22 ;
      RECT 145.22 305.04 149.93 305.2 ;
      RECT 7.38 303.99 88.22 304.33 ;
      RECT 144.57 304.08 149.93 304.24 ;
      RECT 145.22 303.12 149.93 303.28 ;
      RECT 6.24 302.06 7.14 302.86 ;
      RECT 149.63 302.1 149.93 302.8 ;
      RECT 145.22 301.64 149.93 301.8 ;
      RECT 7.38 300.59 88.22 300.93 ;
      RECT 144.63 300.68 149.93 300.84 ;
      RECT 145.22 299.72 149.93 299.88 ;
      RECT 6.24 298.66 7.14 299.46 ;
      RECT 149.63 298.72 149.93 299.42 ;
      RECT 145.22 298.24 149.93 298.4 ;
      RECT 7.38 297.19 88.22 297.53 ;
      RECT 144.57 297.28 149.93 297.44 ;
      RECT 145.22 296.32 149.93 296.48 ;
      RECT 6.24 295.26 7.14 296.06 ;
      RECT 149.63 295.3 149.93 296 ;
      RECT 145.22 294.84 149.93 295 ;
      RECT 7.38 293.79 88.22 294.13 ;
      RECT 144.63 293.88 149.93 294.04 ;
      RECT 145.22 292.92 149.93 293.08 ;
      RECT 6.24 291.86 7.14 292.66 ;
      RECT 149.63 291.92 149.93 292.62 ;
      RECT 145.22 291.44 149.93 291.6 ;
      RECT 7.38 290.39 88.22 290.73 ;
      RECT 144.57 290.48 149.93 290.64 ;
      RECT 145.22 289.52 149.93 289.68 ;
      RECT 6.24 288.46 7.14 289.26 ;
      RECT 149.63 288.5 149.93 289.2 ;
      RECT 145.22 288.04 149.93 288.2 ;
      RECT 7.38 286.99 88.22 287.33 ;
      RECT 144.63 287.08 149.93 287.24 ;
      RECT 145.22 286.12 149.93 286.28 ;
      RECT 6.24 285.06 7.14 285.86 ;
      RECT 149.63 285.12 149.93 285.82 ;
      RECT 145.22 284.64 149.93 284.8 ;
      RECT 7.38 283.59 88.22 283.93 ;
      RECT 144.57 283.68 149.93 283.84 ;
      RECT 145.22 282.72 149.93 282.88 ;
      RECT 6.24 281.66 7.14 282.46 ;
      RECT 149.63 281.7 149.93 282.4 ;
      RECT 145.22 281.24 149.93 281.4 ;
      RECT 7.38 280.19 88.22 280.53 ;
      RECT 144.63 280.28 149.93 280.44 ;
      RECT 145.22 279.32 149.93 279.48 ;
      RECT 6.24 278.26 7.14 279.06 ;
      RECT 149.63 278.32 149.93 279.02 ;
      RECT 145.22 277.84 149.93 278 ;
      RECT 7.38 276.79 88.22 277.13 ;
      RECT 144.57 276.88 149.93 277.04 ;
      RECT 145.22 275.92 149.93 276.08 ;
      RECT 6.24 274.86 7.14 275.66 ;
      RECT 149.63 274.9 149.93 275.6 ;
      RECT 145.22 274.44 149.93 274.6 ;
      RECT 7.38 273.39 88.22 273.73 ;
      RECT 144.63 273.48 149.93 273.64 ;
      RECT 145.22 272.52 149.93 272.68 ;
      RECT 6.24 271.46 7.14 272.26 ;
      RECT 149.63 271.52 149.93 272.22 ;
      RECT 145.22 271.04 149.93 271.2 ;
      RECT 7.38 269.99 88.22 270.33 ;
      RECT 144.57 270.08 149.93 270.24 ;
      RECT 145.22 269.12 149.93 269.28 ;
      RECT 6.24 268.06 7.14 268.86 ;
      RECT 149.63 268.1 149.93 268.8 ;
      RECT 145.22 267.64 149.93 267.8 ;
      RECT 7.38 266.59 88.22 266.93 ;
      RECT 144.63 266.68 149.93 266.84 ;
      RECT 145.22 265.72 149.93 265.88 ;
      RECT 6.24 264.66 7.14 265.46 ;
      RECT 149.63 264.72 149.93 265.42 ;
      RECT 145.22 264.24 149.93 264.4 ;
      RECT 7.38 263.19 88.22 263.53 ;
      RECT 144.57 263.28 149.93 263.44 ;
      RECT 145.22 262.32 149.93 262.48 ;
      RECT 6.24 261.26 7.14 262.06 ;
      RECT 149.63 261.3 149.93 262 ;
      RECT 145.22 260.84 149.93 261 ;
      RECT 7.38 259.79 88.22 260.13 ;
      RECT 144.63 259.88 149.93 260.04 ;
      RECT 145.22 258.92 149.93 259.08 ;
      RECT 6.24 257.86 7.14 258.66 ;
      RECT 149.63 257.92 149.93 258.62 ;
      RECT 145.22 257.44 149.93 257.6 ;
      RECT 7.38 256.39 88.22 256.73 ;
      RECT 144.57 256.48 149.93 256.64 ;
      RECT 145.22 255.52 149.93 255.68 ;
      RECT 6.24 254.46 7.14 255.26 ;
      RECT 149.63 254.5 149.93 255.2 ;
      RECT 145.22 254.04 149.93 254.2 ;
      RECT 7.38 252.99 88.22 253.33 ;
      RECT 144.63 253.08 149.93 253.24 ;
      RECT 145.22 252.12 149.93 252.28 ;
      RECT 6.24 251.06 7.14 251.86 ;
      RECT 149.63 251.12 149.93 251.82 ;
      RECT 145.22 250.64 149.93 250.8 ;
      RECT 7.38 249.59 88.22 249.93 ;
      RECT 144.57 249.68 149.93 249.84 ;
      RECT 145.22 248.72 149.93 248.88 ;
      RECT 6.24 247.66 7.14 248.46 ;
      RECT 149.63 247.7 149.93 248.4 ;
      RECT 145.22 247.24 149.93 247.4 ;
      RECT 7.38 246.19 88.22 246.53 ;
      RECT 144.63 246.28 149.93 246.44 ;
      RECT 145.22 245.32 149.93 245.48 ;
      RECT 6.24 244.26 7.14 245.06 ;
      RECT 149.63 244.32 149.93 245.02 ;
      RECT 145.22 243.84 149.93 244 ;
      RECT 7.38 242.79 88.22 243.13 ;
      RECT 144.57 242.88 149.93 243.04 ;
      RECT 145.22 241.92 149.93 242.08 ;
      RECT 6.24 240.86 7.14 241.66 ;
      RECT 149.63 240.9 149.93 241.6 ;
      RECT 145.22 240.44 149.93 240.6 ;
      RECT 7.38 239.39 88.22 239.73 ;
      RECT 144.63 239.48 149.93 239.64 ;
      RECT 145.22 238.52 149.93 238.68 ;
      RECT 6.24 237.46 7.14 238.26 ;
      RECT 149.63 237.52 149.93 238.22 ;
      RECT 145.22 237.04 149.93 237.2 ;
      RECT 7.38 235.99 88.22 236.33 ;
      RECT 144.57 236.08 149.93 236.24 ;
      RECT 145.22 235.12 149.93 235.28 ;
      RECT 6.24 234.06 7.14 234.86 ;
      RECT 149.63 234.1 149.93 234.8 ;
      RECT 145.22 233.64 149.93 233.8 ;
      RECT 7.38 232.59 88.22 232.93 ;
      RECT 144.63 232.68 149.93 232.84 ;
      RECT 145.22 231.72 149.93 231.88 ;
      RECT 6.24 230.66 7.14 231.46 ;
      RECT 149.63 230.72 149.93 231.42 ;
      RECT 145.22 230.24 149.93 230.4 ;
      RECT 7.38 229.19 88.22 229.53 ;
      RECT 144.57 229.28 149.93 229.44 ;
      RECT 145.22 228.32 149.93 228.48 ;
      RECT 6.24 227.26 7.14 228.06 ;
      RECT 149.63 227.3 149.93 228 ;
      RECT 145.22 226.84 149.93 227 ;
      RECT 7.38 225.79 88.22 226.13 ;
      RECT 144.63 225.88 149.93 226.04 ;
      RECT 145.22 224.92 149.93 225.08 ;
      RECT 6.24 223.86 7.14 224.66 ;
      RECT 149.63 223.92 149.93 224.62 ;
      RECT 145.22 223.44 149.93 223.6 ;
      RECT 7.38 222.39 88.22 222.73 ;
      RECT 144.57 222.48 149.93 222.64 ;
      RECT 145.22 221.52 149.93 221.68 ;
      RECT 6.24 220.46 7.14 221.26 ;
      RECT 149.63 220.5 149.93 221.2 ;
      RECT 145.22 220.04 149.93 220.2 ;
      RECT 7.38 218.99 88.22 219.33 ;
      RECT 144.63 219.08 149.93 219.24 ;
      RECT 145.22 218.12 149.93 218.28 ;
      RECT 6.24 217.06 7.14 217.86 ;
      RECT 149.63 217.12 149.93 217.82 ;
      RECT 145.22 216.64 149.93 216.8 ;
      RECT 7.38 215.59 88.22 215.93 ;
      RECT 144.57 215.68 149.93 215.84 ;
      RECT 145.22 214.72 149.93 214.88 ;
      RECT 6.24 213.66 7.14 214.46 ;
      RECT 149.63 213.7 149.93 214.4 ;
      RECT 145.22 213.24 149.93 213.4 ;
      RECT 7.38 212.19 88.22 212.53 ;
      RECT 144.63 212.28 149.93 212.44 ;
      RECT 145.22 211.32 149.93 211.48 ;
      RECT 6.24 210.26 7.14 211.06 ;
      RECT 149.63 210.32 149.93 211.02 ;
      RECT 145.22 209.84 149.93 210 ;
      RECT 7.38 208.79 88.22 209.13 ;
      RECT 144.57 208.88 149.93 209.04 ;
      RECT 145.22 207.92 149.93 208.08 ;
      RECT 6.24 206.86 7.14 207.66 ;
      RECT 149.63 206.9 149.93 207.6 ;
      RECT 145.22 206.44 149.93 206.6 ;
      RECT 7.38 205.39 88.22 205.73 ;
      RECT 144.63 205.48 149.93 205.64 ;
      RECT 145.22 204.52 149.93 204.68 ;
      RECT 6.24 203.46 7.14 204.26 ;
      RECT 149.63 203.52 149.93 204.22 ;
      RECT 145.22 203.04 149.93 203.2 ;
      RECT 7.38 201.99 88.22 202.33 ;
      RECT 144.57 202.08 149.93 202.24 ;
      RECT 145.22 201.12 149.93 201.28 ;
      RECT 6.24 200.06 7.14 200.86 ;
      RECT 149.63 200.1 149.93 200.8 ;
      RECT 145.22 199.64 149.93 199.8 ;
      RECT 7.38 198.59 88.22 198.93 ;
      RECT 144.63 198.68 149.93 198.84 ;
      RECT 145.22 197.72 149.93 197.88 ;
      RECT 6.24 196.66 7.14 197.46 ;
      RECT 149.63 196.72 149.93 197.42 ;
      RECT 145.22 196.24 149.93 196.4 ;
      RECT 7.38 195.19 88.22 195.53 ;
      RECT 144.57 195.28 149.93 195.44 ;
      RECT 145.22 194.32 149.93 194.48 ;
      RECT 6.24 193.26 7.14 194.06 ;
      RECT 149.63 193.3 149.93 194 ;
      RECT 145.22 192.84 149.93 193 ;
      RECT 7.38 191.79 88.22 192.13 ;
      RECT 144.63 191.88 149.93 192.04 ;
      RECT 145.22 190.92 149.93 191.08 ;
      RECT 6.24 189.86 7.14 190.66 ;
      RECT 149.63 189.92 149.93 190.62 ;
      RECT 145.22 189.44 149.93 189.6 ;
      RECT 7.38 188.39 88.22 188.73 ;
      RECT 144.57 188.48 149.93 188.64 ;
      RECT 145.22 187.52 149.93 187.68 ;
      RECT 6.24 186.46 7.14 187.26 ;
      RECT 149.63 186.5 149.93 187.2 ;
      RECT 145.22 186.04 149.93 186.2 ;
      RECT 7.38 184.99 88.22 185.33 ;
      RECT 144.63 185.08 149.93 185.24 ;
      RECT 145.22 184.12 149.93 184.28 ;
      RECT 6.24 183.06 7.14 183.86 ;
      RECT 149.63 183.12 149.93 183.82 ;
      RECT 145.22 182.64 149.93 182.8 ;
      RECT 7.38 181.59 88.22 181.93 ;
      RECT 144.57 181.68 149.93 181.84 ;
      RECT 145.22 180.72 149.93 180.88 ;
      RECT 6.24 179.66 7.14 180.46 ;
      RECT 149.63 179.7 149.93 180.4 ;
      RECT 145.22 179.24 149.93 179.4 ;
      RECT 7.38 178.19 88.22 178.53 ;
      RECT 144.63 178.28 149.93 178.44 ;
      RECT 145.22 177.32 149.93 177.48 ;
      RECT 6.24 176.26 7.14 177.06 ;
      RECT 149.63 176.32 149.93 177.02 ;
      RECT 145.22 175.84 149.93 176 ;
      RECT 7.38 174.79 88.22 175.13 ;
      RECT 144.57 174.88 149.93 175.04 ;
      RECT 145.22 173.92 149.93 174.08 ;
      RECT 6.24 172.86 7.14 173.66 ;
      RECT 149.63 172.9 149.93 173.6 ;
      RECT 145.22 172.44 149.93 172.6 ;
      RECT 7.38 171.39 88.22 171.73 ;
      RECT 144.63 171.48 149.93 171.64 ;
      RECT 145.22 170.52 149.93 170.68 ;
      RECT 6.24 169.46 7.14 170.26 ;
      RECT 149.63 169.52 149.93 170.22 ;
      RECT 145.22 169.04 149.93 169.2 ;
      RECT 7.38 167.99 88.22 168.33 ;
      RECT 144.57 168.08 149.93 168.24 ;
      RECT 145.22 167.12 149.93 167.28 ;
      RECT 6.24 166.06 7.14 166.86 ;
      RECT 149.63 166.1 149.93 166.8 ;
      RECT 145.22 165.64 149.93 165.8 ;
      RECT 7.38 164.59 88.22 164.93 ;
      RECT 144.63 164.68 149.93 164.84 ;
      RECT 145.22 163.72 149.93 163.88 ;
      RECT 6.24 162.66 7.14 163.46 ;
      RECT 149.63 162.72 149.93 163.42 ;
      RECT 145.22 162.24 149.93 162.4 ;
      RECT 7.38 161.19 88.22 161.53 ;
      RECT 144.57 161.28 149.93 161.44 ;
      RECT 145.22 160.32 149.93 160.48 ;
      RECT 6.24 159.26 7.14 160.06 ;
      RECT 149.63 159.3 149.93 160 ;
      RECT 145.22 158.84 149.93 159 ;
      RECT 7.38 157.79 88.22 158.13 ;
      RECT 144.63 157.88 149.93 158.04 ;
      RECT 145.22 156.92 149.93 157.08 ;
      RECT 6.24 155.86 7.14 156.66 ;
      RECT 149.63 155.92 149.93 156.62 ;
      RECT 145.22 155.44 149.93 155.6 ;
      RECT 7.38 154.39 88.22 154.73 ;
      RECT 144.57 154.48 149.93 154.64 ;
      RECT 6.24 152.46 7.14 153.26 ;
      RECT 7.38 150.99 88.22 151.33 ;
      RECT 6.24 149.06 7.14 149.86 ;
      RECT 7.38 147.59 88.22 147.93 ;
      RECT 6.24 145.66 7.14 146.46 ;
      RECT 7.38 144.19 88.22 144.53 ;
      RECT 6.24 142.26 7.14 143.06 ;
      RECT 7.38 140.79 88.22 141.13 ;
      RECT 6.24 138.86 7.14 139.66 ;
      RECT 7.38 137.39 88.22 137.73 ;
      RECT 6.24 135.46 7.14 136.26 ;
      RECT 7.38 133.99 88.22 134.33 ;
      RECT 6.24 132.06 7.14 132.86 ;
      RECT 7.38 130.59 88.22 130.93 ;
      RECT 6.24 128.66 7.14 129.46 ;
      RECT 7.38 127.19 88.22 127.53 ;
      RECT 6.24 125.26 7.14 126.06 ;
      RECT 7.38 123.79 88.22 124.13 ;
      RECT 6.24 121.86 7.14 122.66 ;
      RECT 7.38 120.39 88.22 120.73 ;
      RECT 6.24 118.46 7.14 119.26 ;
      RECT 7.38 116.99 88.22 117.33 ;
      RECT 6.24 115.06 7.14 115.86 ;
      RECT 7.38 113.59 88.22 113.93 ;
      RECT 6.24 111.66 7.14 112.46 ;
      RECT 7.38 110.19 88.22 110.53 ;
      RECT 6.24 108.26 7.14 109.06 ;
      RECT 7.38 106.79 88.22 107.13 ;
      RECT 6.24 104.86 7.14 105.66 ;
      RECT 7.38 103.39 88.22 103.73 ;
      RECT 6.24 101.46 7.14 102.26 ;
      RECT 7.38 99.99 88.22 100.33 ;
      RECT 6.24 98.06 7.14 98.86 ;
      RECT 7.38 96.59 88.22 96.93 ;
      RECT 6.24 94.66 7.14 95.46 ;
      RECT 7.38 93.19 88.22 93.53 ;
      RECT 6.24 91.26 7.14 92.06 ;
      RECT 7.38 89.79 88.22 90.13 ;
      RECT 6.24 87.86 7.14 88.66 ;
      RECT 7.38 86.39 88.22 86.73 ;
      RECT 6.24 84.46 7.14 85.26 ;
      RECT 7.38 82.99 88.22 83.33 ;
      RECT 6.24 81.06 7.14 81.86 ;
      RECT 7.38 79.59 88.22 79.93 ;
      RECT 6.24 77.66 7.14 78.46 ;
      RECT 7.38 76.19 88.22 76.53 ;
      RECT 6.24 74.26 7.14 75.06 ;
      RECT 7.38 72.79 88.22 73.13 ;
      RECT 6.24 70.86 7.14 71.66 ;
      RECT 7.38 69.46 88.22 69.73 ;
      RECT 6.98 69.07 87.44 69.3 ;
      RECT 86.8 67.1 87 509.88 ;
      RECT 6.98 67.81 7.46 68.09 ;
      RECT 7.24 8.2 7.46 68.09 ;
      RECT 86.8 67.1 87.9 67.3 ;
      RECT 87.62 21.41 87.9 67.3 ;
      RECT 6.24 54.22 7.46 55.22 ;
      RECT 6.24 41.29 7.46 42.29 ;
      RECT 6.24 39.44 7.46 40.44 ;
      RECT 6.24 32.98 7.46 33.98 ;
      RECT 6.24 31.13 7.46 32.13 ;
      RECT 6.24 21.41 7.46 22.21 ;
      RECT 6.24 12.64 7.46 13.74 ;
      RECT 147.93 30.63 148.09 32.23 ;
      RECT 147.93 30.63 148.27 30.79 ;
      RECT 148.11 29.46 148.27 30.79 ;
      RECT 147.61 29.46 149.63 29.62 ;
      RECT 147.61 27.81 147.77 29.62 ;
      RECT 148.05 509.72 149.61 509.88 ;
      RECT 149.45 506.88 149.61 509.88 ;
      RECT 148.73 506.88 149.61 507.04 ;
      RECT 149.39 30.1 149.55 32.94 ;
      RECT 149.39 32.26 149.56 32.58 ;
      RECT 149.17 30.1 149.55 30.26 ;
      RECT 143.1 71 145.06 71.16 ;
      RECT 144.8 69.96 145.06 71.16 ;
      RECT 144.8 70.92 149.4 71.08 ;
      RECT 135.8 70.92 143.38 71.08 ;
      RECT 135.8 69.96 149.4 70.12 ;
      RECT 135.8 72.4 149.4 72.56 ;
      RECT 144.8 71.36 145.06 72.56 ;
      RECT 144.8 71.44 149.4 71.6 ;
      RECT 135.8 71.44 143.38 71.6 ;
      RECT 143.1 71.36 145.06 71.52 ;
      RECT 143.1 74.4 145.06 74.56 ;
      RECT 144.8 73.36 145.06 74.56 ;
      RECT 144.8 74.32 149.4 74.48 ;
      RECT 135.8 74.32 143.38 74.48 ;
      RECT 135.8 73.36 149.4 73.52 ;
      RECT 135.8 75.8 149.4 75.96 ;
      RECT 144.8 74.76 145.06 75.96 ;
      RECT 144.8 74.84 149.4 75 ;
      RECT 135.8 74.84 143.38 75 ;
      RECT 143.1 74.76 145.06 74.92 ;
      RECT 143.1 77.8 145.06 77.96 ;
      RECT 144.8 76.76 145.06 77.96 ;
      RECT 144.8 77.72 149.4 77.88 ;
      RECT 135.8 77.72 143.38 77.88 ;
      RECT 135.8 76.76 149.4 76.92 ;
      RECT 135.8 79.2 149.4 79.36 ;
      RECT 144.8 78.16 145.06 79.36 ;
      RECT 144.8 78.24 149.4 78.4 ;
      RECT 135.8 78.24 143.38 78.4 ;
      RECT 143.1 78.16 145.06 78.32 ;
      RECT 143.1 81.2 145.06 81.36 ;
      RECT 144.8 80.16 145.06 81.36 ;
      RECT 144.8 81.12 149.4 81.28 ;
      RECT 135.8 81.12 143.38 81.28 ;
      RECT 135.8 80.16 149.4 80.32 ;
      RECT 135.8 82.6 149.4 82.76 ;
      RECT 144.8 81.56 145.06 82.76 ;
      RECT 144.8 81.64 149.4 81.8 ;
      RECT 135.8 81.64 143.38 81.8 ;
      RECT 143.1 81.56 145.06 81.72 ;
      RECT 143.1 84.6 145.06 84.76 ;
      RECT 144.8 83.56 145.06 84.76 ;
      RECT 144.8 84.52 149.4 84.68 ;
      RECT 135.8 84.52 143.38 84.68 ;
      RECT 135.8 83.56 149.4 83.72 ;
      RECT 135.8 86 149.4 86.16 ;
      RECT 144.8 84.96 145.06 86.16 ;
      RECT 144.8 85.04 149.4 85.2 ;
      RECT 135.8 85.04 143.38 85.2 ;
      RECT 143.1 84.96 145.06 85.12 ;
      RECT 143.1 88 145.06 88.16 ;
      RECT 144.8 86.96 145.06 88.16 ;
      RECT 144.8 87.92 149.4 88.08 ;
      RECT 135.8 87.92 143.38 88.08 ;
      RECT 135.8 86.96 149.4 87.12 ;
      RECT 135.8 89.4 149.4 89.56 ;
      RECT 144.8 88.36 145.06 89.56 ;
      RECT 144.8 88.44 149.4 88.6 ;
      RECT 135.8 88.44 143.38 88.6 ;
      RECT 143.1 88.36 145.06 88.52 ;
      RECT 143.1 91.4 145.06 91.56 ;
      RECT 144.8 90.36 145.06 91.56 ;
      RECT 144.8 91.32 149.4 91.48 ;
      RECT 135.8 91.32 143.38 91.48 ;
      RECT 135.8 90.36 149.4 90.52 ;
      RECT 135.8 92.8 149.4 92.96 ;
      RECT 144.8 91.76 145.06 92.96 ;
      RECT 144.8 91.84 149.4 92 ;
      RECT 135.8 91.84 143.38 92 ;
      RECT 143.1 91.76 145.06 91.92 ;
      RECT 143.1 94.8 145.06 94.96 ;
      RECT 144.8 93.76 145.06 94.96 ;
      RECT 144.8 94.72 149.4 94.88 ;
      RECT 135.8 94.72 143.38 94.88 ;
      RECT 135.8 93.76 149.4 93.92 ;
      RECT 135.8 96.2 149.4 96.36 ;
      RECT 144.8 95.16 145.06 96.36 ;
      RECT 144.8 95.24 149.4 95.4 ;
      RECT 135.8 95.24 143.38 95.4 ;
      RECT 143.1 95.16 145.06 95.32 ;
      RECT 143.1 98.2 145.06 98.36 ;
      RECT 144.8 97.16 145.06 98.36 ;
      RECT 144.8 98.12 149.4 98.28 ;
      RECT 135.8 98.12 143.38 98.28 ;
      RECT 135.8 97.16 149.4 97.32 ;
      RECT 135.8 99.6 149.4 99.76 ;
      RECT 144.8 98.56 145.06 99.76 ;
      RECT 144.8 98.64 149.4 98.8 ;
      RECT 135.8 98.64 143.38 98.8 ;
      RECT 143.1 98.56 145.06 98.72 ;
      RECT 143.1 101.6 145.06 101.76 ;
      RECT 144.8 100.56 145.06 101.76 ;
      RECT 144.8 101.52 149.4 101.68 ;
      RECT 135.8 101.52 143.38 101.68 ;
      RECT 135.8 100.56 149.4 100.72 ;
      RECT 135.8 103 149.4 103.16 ;
      RECT 144.8 101.96 145.06 103.16 ;
      RECT 144.8 102.04 149.4 102.2 ;
      RECT 135.8 102.04 143.38 102.2 ;
      RECT 143.1 101.96 145.06 102.12 ;
      RECT 143.1 105 145.06 105.16 ;
      RECT 144.8 103.96 145.06 105.16 ;
      RECT 144.8 104.92 149.4 105.08 ;
      RECT 135.8 104.92 143.38 105.08 ;
      RECT 135.8 103.96 149.4 104.12 ;
      RECT 135.8 106.4 149.4 106.56 ;
      RECT 144.8 105.36 145.06 106.56 ;
      RECT 144.8 105.44 149.4 105.6 ;
      RECT 135.8 105.44 143.38 105.6 ;
      RECT 143.1 105.36 145.06 105.52 ;
      RECT 143.1 108.4 145.06 108.56 ;
      RECT 144.8 107.36 145.06 108.56 ;
      RECT 144.8 108.32 149.4 108.48 ;
      RECT 135.8 108.32 143.38 108.48 ;
      RECT 135.8 107.36 149.4 107.52 ;
      RECT 135.8 109.8 149.4 109.96 ;
      RECT 144.8 108.76 145.06 109.96 ;
      RECT 144.8 108.84 149.4 109 ;
      RECT 135.8 108.84 143.38 109 ;
      RECT 143.1 108.76 145.06 108.92 ;
      RECT 143.1 111.8 145.06 111.96 ;
      RECT 144.8 110.76 145.06 111.96 ;
      RECT 144.8 111.72 149.4 111.88 ;
      RECT 135.8 111.72 143.38 111.88 ;
      RECT 135.8 110.76 149.4 110.92 ;
      RECT 135.8 113.2 149.4 113.36 ;
      RECT 144.8 112.16 145.06 113.36 ;
      RECT 144.8 112.24 149.4 112.4 ;
      RECT 135.8 112.24 143.38 112.4 ;
      RECT 143.1 112.16 145.06 112.32 ;
      RECT 143.1 115.2 145.06 115.36 ;
      RECT 144.8 114.16 145.06 115.36 ;
      RECT 144.8 115.12 149.4 115.28 ;
      RECT 135.8 115.12 143.38 115.28 ;
      RECT 135.8 114.16 149.4 114.32 ;
      RECT 135.8 116.6 149.4 116.76 ;
      RECT 144.8 115.56 145.06 116.76 ;
      RECT 144.8 115.64 149.4 115.8 ;
      RECT 135.8 115.64 143.38 115.8 ;
      RECT 143.1 115.56 145.06 115.72 ;
      RECT 143.1 118.6 145.06 118.76 ;
      RECT 144.8 117.56 145.06 118.76 ;
      RECT 144.8 118.52 149.4 118.68 ;
      RECT 135.8 118.52 143.38 118.68 ;
      RECT 135.8 117.56 149.4 117.72 ;
      RECT 135.8 120 149.4 120.16 ;
      RECT 144.8 118.96 145.06 120.16 ;
      RECT 144.8 119.04 149.4 119.2 ;
      RECT 135.8 119.04 143.38 119.2 ;
      RECT 143.1 118.96 145.06 119.12 ;
      RECT 143.1 122 145.06 122.16 ;
      RECT 144.8 120.96 145.06 122.16 ;
      RECT 144.8 121.92 149.4 122.08 ;
      RECT 135.8 121.92 143.38 122.08 ;
      RECT 135.8 120.96 149.4 121.12 ;
      RECT 135.8 123.4 149.4 123.56 ;
      RECT 144.8 122.36 145.06 123.56 ;
      RECT 144.8 122.44 149.4 122.6 ;
      RECT 135.8 122.44 143.38 122.6 ;
      RECT 143.1 122.36 145.06 122.52 ;
      RECT 143.1 125.4 145.06 125.56 ;
      RECT 144.8 124.36 145.06 125.56 ;
      RECT 144.8 125.32 149.4 125.48 ;
      RECT 135.8 125.32 143.38 125.48 ;
      RECT 135.8 124.36 149.4 124.52 ;
      RECT 135.8 126.8 149.4 126.96 ;
      RECT 144.8 125.76 145.06 126.96 ;
      RECT 144.8 125.84 149.4 126 ;
      RECT 135.8 125.84 143.38 126 ;
      RECT 143.1 125.76 145.06 125.92 ;
      RECT 143.1 128.8 145.06 128.96 ;
      RECT 144.8 127.76 145.06 128.96 ;
      RECT 144.8 128.72 149.4 128.88 ;
      RECT 135.8 128.72 143.38 128.88 ;
      RECT 135.8 127.76 149.4 127.92 ;
      RECT 135.8 130.2 149.4 130.36 ;
      RECT 144.8 129.16 145.06 130.36 ;
      RECT 144.8 129.24 149.4 129.4 ;
      RECT 135.8 129.24 143.38 129.4 ;
      RECT 143.1 129.16 145.06 129.32 ;
      RECT 143.1 132.2 145.06 132.36 ;
      RECT 144.8 131.16 145.06 132.36 ;
      RECT 144.8 132.12 149.4 132.28 ;
      RECT 135.8 132.12 143.38 132.28 ;
      RECT 135.8 131.16 149.4 131.32 ;
      RECT 135.8 133.6 149.4 133.76 ;
      RECT 144.8 132.56 145.06 133.76 ;
      RECT 144.8 132.64 149.4 132.8 ;
      RECT 135.8 132.64 143.38 132.8 ;
      RECT 143.1 132.56 145.06 132.72 ;
      RECT 143.1 135.6 145.06 135.76 ;
      RECT 144.8 134.56 145.06 135.76 ;
      RECT 144.8 135.52 149.4 135.68 ;
      RECT 135.8 135.52 143.38 135.68 ;
      RECT 135.8 134.56 149.4 134.72 ;
      RECT 135.8 137 149.4 137.16 ;
      RECT 144.8 135.96 145.06 137.16 ;
      RECT 144.8 136.04 149.4 136.2 ;
      RECT 135.8 136.04 143.38 136.2 ;
      RECT 143.1 135.96 145.06 136.12 ;
      RECT 143.1 139 145.06 139.16 ;
      RECT 144.8 137.96 145.06 139.16 ;
      RECT 144.8 138.92 149.4 139.08 ;
      RECT 135.8 138.92 143.38 139.08 ;
      RECT 135.8 137.96 149.4 138.12 ;
      RECT 135.8 140.4 149.4 140.56 ;
      RECT 144.8 139.36 145.06 140.56 ;
      RECT 144.8 139.44 149.4 139.6 ;
      RECT 135.8 139.44 143.38 139.6 ;
      RECT 143.1 139.36 145.06 139.52 ;
      RECT 143.1 142.4 145.06 142.56 ;
      RECT 144.8 141.36 145.06 142.56 ;
      RECT 144.8 142.32 149.4 142.48 ;
      RECT 135.8 142.32 143.38 142.48 ;
      RECT 135.8 141.36 149.4 141.52 ;
      RECT 135.8 143.8 149.4 143.96 ;
      RECT 144.8 142.76 145.06 143.96 ;
      RECT 144.8 142.84 149.4 143 ;
      RECT 135.8 142.84 143.38 143 ;
      RECT 143.1 142.76 145.06 142.92 ;
      RECT 143.1 145.8 145.06 145.96 ;
      RECT 144.8 144.76 145.06 145.96 ;
      RECT 144.8 145.72 149.4 145.88 ;
      RECT 135.8 145.72 143.38 145.88 ;
      RECT 135.8 144.76 149.4 144.92 ;
      RECT 135.8 147.2 149.4 147.36 ;
      RECT 144.8 146.16 145.06 147.36 ;
      RECT 144.8 146.24 149.4 146.4 ;
      RECT 135.8 146.24 143.38 146.4 ;
      RECT 143.1 146.16 145.06 146.32 ;
      RECT 143.1 149.2 145.06 149.36 ;
      RECT 144.8 148.16 145.06 149.36 ;
      RECT 144.8 149.12 149.4 149.28 ;
      RECT 135.8 149.12 143.38 149.28 ;
      RECT 135.8 148.16 149.4 148.32 ;
      RECT 135.8 150.6 149.4 150.76 ;
      RECT 144.8 149.56 145.06 150.76 ;
      RECT 144.8 149.64 149.4 149.8 ;
      RECT 135.8 149.64 143.38 149.8 ;
      RECT 143.1 149.56 145.06 149.72 ;
      RECT 143.1 152.6 145.06 152.76 ;
      RECT 144.8 151.56 145.06 152.76 ;
      RECT 144.8 152.52 149.4 152.68 ;
      RECT 135.8 152.52 143.38 152.68 ;
      RECT 135.8 151.56 149.4 151.72 ;
      RECT 135.8 154 149.4 154.16 ;
      RECT 144.8 152.96 145.06 154.16 ;
      RECT 144.8 153.04 149.4 153.2 ;
      RECT 135.8 153.04 143.38 153.2 ;
      RECT 143.1 152.96 145.06 153.12 ;
      RECT 143.1 156 145.06 156.16 ;
      RECT 144.8 154.96 145.06 156.16 ;
      RECT 144.8 155.92 149.4 156.08 ;
      RECT 135.8 155.92 143.38 156.08 ;
      RECT 135.8 154.96 149.4 155.12 ;
      RECT 135.8 157.4 149.4 157.56 ;
      RECT 144.8 156.36 145.06 157.56 ;
      RECT 144.8 156.44 149.4 156.6 ;
      RECT 135.8 156.44 143.38 156.6 ;
      RECT 143.1 156.36 145.06 156.52 ;
      RECT 143.1 159.4 145.06 159.56 ;
      RECT 144.8 158.36 145.06 159.56 ;
      RECT 144.8 159.32 149.4 159.48 ;
      RECT 135.8 159.32 143.38 159.48 ;
      RECT 135.8 158.36 149.4 158.52 ;
      RECT 135.8 160.8 149.4 160.96 ;
      RECT 144.8 159.76 145.06 160.96 ;
      RECT 144.8 159.84 149.4 160 ;
      RECT 135.8 159.84 143.38 160 ;
      RECT 143.1 159.76 145.06 159.92 ;
      RECT 143.1 162.8 145.06 162.96 ;
      RECT 144.8 161.76 145.06 162.96 ;
      RECT 144.8 162.72 149.4 162.88 ;
      RECT 135.8 162.72 143.38 162.88 ;
      RECT 135.8 161.76 149.4 161.92 ;
      RECT 135.8 164.2 149.4 164.36 ;
      RECT 144.8 163.16 145.06 164.36 ;
      RECT 144.8 163.24 149.4 163.4 ;
      RECT 135.8 163.24 143.38 163.4 ;
      RECT 143.1 163.16 145.06 163.32 ;
      RECT 143.1 166.2 145.06 166.36 ;
      RECT 144.8 165.16 145.06 166.36 ;
      RECT 144.8 166.12 149.4 166.28 ;
      RECT 135.8 166.12 143.38 166.28 ;
      RECT 135.8 165.16 149.4 165.32 ;
      RECT 135.8 167.6 149.4 167.76 ;
      RECT 144.8 166.56 145.06 167.76 ;
      RECT 144.8 166.64 149.4 166.8 ;
      RECT 135.8 166.64 143.38 166.8 ;
      RECT 143.1 166.56 145.06 166.72 ;
      RECT 143.1 169.6 145.06 169.76 ;
      RECT 144.8 168.56 145.06 169.76 ;
      RECT 144.8 169.52 149.4 169.68 ;
      RECT 135.8 169.52 143.38 169.68 ;
      RECT 135.8 168.56 149.4 168.72 ;
      RECT 135.8 171 149.4 171.16 ;
      RECT 144.8 169.96 145.06 171.16 ;
      RECT 144.8 170.04 149.4 170.2 ;
      RECT 135.8 170.04 143.38 170.2 ;
      RECT 143.1 169.96 145.06 170.12 ;
      RECT 143.1 173 145.06 173.16 ;
      RECT 144.8 171.96 145.06 173.16 ;
      RECT 144.8 172.92 149.4 173.08 ;
      RECT 135.8 172.92 143.38 173.08 ;
      RECT 135.8 171.96 149.4 172.12 ;
      RECT 135.8 174.4 149.4 174.56 ;
      RECT 144.8 173.36 145.06 174.56 ;
      RECT 144.8 173.44 149.4 173.6 ;
      RECT 135.8 173.44 143.38 173.6 ;
      RECT 143.1 173.36 145.06 173.52 ;
      RECT 143.1 176.4 145.06 176.56 ;
      RECT 144.8 175.36 145.06 176.56 ;
      RECT 144.8 176.32 149.4 176.48 ;
      RECT 135.8 176.32 143.38 176.48 ;
      RECT 135.8 175.36 149.4 175.52 ;
      RECT 135.8 177.8 149.4 177.96 ;
      RECT 144.8 176.76 145.06 177.96 ;
      RECT 144.8 176.84 149.4 177 ;
      RECT 135.8 176.84 143.38 177 ;
      RECT 143.1 176.76 145.06 176.92 ;
      RECT 143.1 179.8 145.06 179.96 ;
      RECT 144.8 178.76 145.06 179.96 ;
      RECT 144.8 179.72 149.4 179.88 ;
      RECT 135.8 179.72 143.38 179.88 ;
      RECT 135.8 178.76 149.4 178.92 ;
      RECT 135.8 181.2 149.4 181.36 ;
      RECT 144.8 180.16 145.06 181.36 ;
      RECT 144.8 180.24 149.4 180.4 ;
      RECT 135.8 180.24 143.38 180.4 ;
      RECT 143.1 180.16 145.06 180.32 ;
      RECT 143.1 183.2 145.06 183.36 ;
      RECT 144.8 182.16 145.06 183.36 ;
      RECT 144.8 183.12 149.4 183.28 ;
      RECT 135.8 183.12 143.38 183.28 ;
      RECT 135.8 182.16 149.4 182.32 ;
      RECT 135.8 184.6 149.4 184.76 ;
      RECT 144.8 183.56 145.06 184.76 ;
      RECT 144.8 183.64 149.4 183.8 ;
      RECT 135.8 183.64 143.38 183.8 ;
      RECT 143.1 183.56 145.06 183.72 ;
      RECT 143.1 186.6 145.06 186.76 ;
      RECT 144.8 185.56 145.06 186.76 ;
      RECT 144.8 186.52 149.4 186.68 ;
      RECT 135.8 186.52 143.38 186.68 ;
      RECT 135.8 185.56 149.4 185.72 ;
      RECT 135.8 188 149.4 188.16 ;
      RECT 144.8 186.96 145.06 188.16 ;
      RECT 144.8 187.04 149.4 187.2 ;
      RECT 135.8 187.04 143.38 187.2 ;
      RECT 143.1 186.96 145.06 187.12 ;
      RECT 143.1 190 145.06 190.16 ;
      RECT 144.8 188.96 145.06 190.16 ;
      RECT 144.8 189.92 149.4 190.08 ;
      RECT 135.8 189.92 143.38 190.08 ;
      RECT 135.8 188.96 149.4 189.12 ;
      RECT 135.8 191.4 149.4 191.56 ;
      RECT 144.8 190.36 145.06 191.56 ;
      RECT 144.8 190.44 149.4 190.6 ;
      RECT 135.8 190.44 143.38 190.6 ;
      RECT 143.1 190.36 145.06 190.52 ;
      RECT 143.1 193.4 145.06 193.56 ;
      RECT 144.8 192.36 145.06 193.56 ;
      RECT 144.8 193.32 149.4 193.48 ;
      RECT 135.8 193.32 143.38 193.48 ;
      RECT 135.8 192.36 149.4 192.52 ;
      RECT 135.8 194.8 149.4 194.96 ;
      RECT 144.8 193.76 145.06 194.96 ;
      RECT 144.8 193.84 149.4 194 ;
      RECT 135.8 193.84 143.38 194 ;
      RECT 143.1 193.76 145.06 193.92 ;
      RECT 143.1 196.8 145.06 196.96 ;
      RECT 144.8 195.76 145.06 196.96 ;
      RECT 144.8 196.72 149.4 196.88 ;
      RECT 135.8 196.72 143.38 196.88 ;
      RECT 135.8 195.76 149.4 195.92 ;
      RECT 135.8 198.2 149.4 198.36 ;
      RECT 144.8 197.16 145.06 198.36 ;
      RECT 144.8 197.24 149.4 197.4 ;
      RECT 135.8 197.24 143.38 197.4 ;
      RECT 143.1 197.16 145.06 197.32 ;
      RECT 143.1 200.2 145.06 200.36 ;
      RECT 144.8 199.16 145.06 200.36 ;
      RECT 144.8 200.12 149.4 200.28 ;
      RECT 135.8 200.12 143.38 200.28 ;
      RECT 135.8 199.16 149.4 199.32 ;
      RECT 135.8 201.6 149.4 201.76 ;
      RECT 144.8 200.56 145.06 201.76 ;
      RECT 144.8 200.64 149.4 200.8 ;
      RECT 135.8 200.64 143.38 200.8 ;
      RECT 143.1 200.56 145.06 200.72 ;
      RECT 143.1 203.6 145.06 203.76 ;
      RECT 144.8 202.56 145.06 203.76 ;
      RECT 144.8 203.52 149.4 203.68 ;
      RECT 135.8 203.52 143.38 203.68 ;
      RECT 135.8 202.56 149.4 202.72 ;
      RECT 135.8 205 149.4 205.16 ;
      RECT 144.8 203.96 145.06 205.16 ;
      RECT 144.8 204.04 149.4 204.2 ;
      RECT 135.8 204.04 143.38 204.2 ;
      RECT 143.1 203.96 145.06 204.12 ;
      RECT 143.1 207 145.06 207.16 ;
      RECT 144.8 205.96 145.06 207.16 ;
      RECT 144.8 206.92 149.4 207.08 ;
      RECT 135.8 206.92 143.38 207.08 ;
      RECT 135.8 205.96 149.4 206.12 ;
      RECT 135.8 208.4 149.4 208.56 ;
      RECT 144.8 207.36 145.06 208.56 ;
      RECT 144.8 207.44 149.4 207.6 ;
      RECT 135.8 207.44 143.38 207.6 ;
      RECT 143.1 207.36 145.06 207.52 ;
      RECT 143.1 210.4 145.06 210.56 ;
      RECT 144.8 209.36 145.06 210.56 ;
      RECT 144.8 210.32 149.4 210.48 ;
      RECT 135.8 210.32 143.38 210.48 ;
      RECT 135.8 209.36 149.4 209.52 ;
      RECT 135.8 211.8 149.4 211.96 ;
      RECT 144.8 210.76 145.06 211.96 ;
      RECT 144.8 210.84 149.4 211 ;
      RECT 135.8 210.84 143.38 211 ;
      RECT 143.1 210.76 145.06 210.92 ;
      RECT 143.1 213.8 145.06 213.96 ;
      RECT 144.8 212.76 145.06 213.96 ;
      RECT 144.8 213.72 149.4 213.88 ;
      RECT 135.8 213.72 143.38 213.88 ;
      RECT 135.8 212.76 149.4 212.92 ;
      RECT 135.8 215.2 149.4 215.36 ;
      RECT 144.8 214.16 145.06 215.36 ;
      RECT 144.8 214.24 149.4 214.4 ;
      RECT 135.8 214.24 143.38 214.4 ;
      RECT 143.1 214.16 145.06 214.32 ;
      RECT 143.1 217.2 145.06 217.36 ;
      RECT 144.8 216.16 145.06 217.36 ;
      RECT 144.8 217.12 149.4 217.28 ;
      RECT 135.8 217.12 143.38 217.28 ;
      RECT 135.8 216.16 149.4 216.32 ;
      RECT 135.8 218.6 149.4 218.76 ;
      RECT 144.8 217.56 145.06 218.76 ;
      RECT 144.8 217.64 149.4 217.8 ;
      RECT 135.8 217.64 143.38 217.8 ;
      RECT 143.1 217.56 145.06 217.72 ;
      RECT 143.1 220.6 145.06 220.76 ;
      RECT 144.8 219.56 145.06 220.76 ;
      RECT 144.8 220.52 149.4 220.68 ;
      RECT 135.8 220.52 143.38 220.68 ;
      RECT 135.8 219.56 149.4 219.72 ;
      RECT 135.8 222 149.4 222.16 ;
      RECT 144.8 220.96 145.06 222.16 ;
      RECT 144.8 221.04 149.4 221.2 ;
      RECT 135.8 221.04 143.38 221.2 ;
      RECT 143.1 220.96 145.06 221.12 ;
      RECT 143.1 224 145.06 224.16 ;
      RECT 144.8 222.96 145.06 224.16 ;
      RECT 144.8 223.92 149.4 224.08 ;
      RECT 135.8 223.92 143.38 224.08 ;
      RECT 135.8 222.96 149.4 223.12 ;
      RECT 135.8 225.4 149.4 225.56 ;
      RECT 144.8 224.36 145.06 225.56 ;
      RECT 144.8 224.44 149.4 224.6 ;
      RECT 135.8 224.44 143.38 224.6 ;
      RECT 143.1 224.36 145.06 224.52 ;
      RECT 143.1 227.4 145.06 227.56 ;
      RECT 144.8 226.36 145.06 227.56 ;
      RECT 144.8 227.32 149.4 227.48 ;
      RECT 135.8 227.32 143.38 227.48 ;
      RECT 135.8 226.36 149.4 226.52 ;
      RECT 135.8 228.8 149.4 228.96 ;
      RECT 144.8 227.76 145.06 228.96 ;
      RECT 144.8 227.84 149.4 228 ;
      RECT 135.8 227.84 143.38 228 ;
      RECT 143.1 227.76 145.06 227.92 ;
      RECT 143.1 230.8 145.06 230.96 ;
      RECT 144.8 229.76 145.06 230.96 ;
      RECT 144.8 230.72 149.4 230.88 ;
      RECT 135.8 230.72 143.38 230.88 ;
      RECT 135.8 229.76 149.4 229.92 ;
      RECT 135.8 232.2 149.4 232.36 ;
      RECT 144.8 231.16 145.06 232.36 ;
      RECT 144.8 231.24 149.4 231.4 ;
      RECT 135.8 231.24 143.38 231.4 ;
      RECT 143.1 231.16 145.06 231.32 ;
      RECT 143.1 234.2 145.06 234.36 ;
      RECT 144.8 233.16 145.06 234.36 ;
      RECT 144.8 234.12 149.4 234.28 ;
      RECT 135.8 234.12 143.38 234.28 ;
      RECT 135.8 233.16 149.4 233.32 ;
      RECT 135.8 235.6 149.4 235.76 ;
      RECT 144.8 234.56 145.06 235.76 ;
      RECT 144.8 234.64 149.4 234.8 ;
      RECT 135.8 234.64 143.38 234.8 ;
      RECT 143.1 234.56 145.06 234.72 ;
      RECT 143.1 237.6 145.06 237.76 ;
      RECT 144.8 236.56 145.06 237.76 ;
      RECT 144.8 237.52 149.4 237.68 ;
      RECT 135.8 237.52 143.38 237.68 ;
      RECT 135.8 236.56 149.4 236.72 ;
      RECT 135.8 239 149.4 239.16 ;
      RECT 144.8 237.96 145.06 239.16 ;
      RECT 144.8 238.04 149.4 238.2 ;
      RECT 135.8 238.04 143.38 238.2 ;
      RECT 143.1 237.96 145.06 238.12 ;
      RECT 143.1 241 145.06 241.16 ;
      RECT 144.8 239.96 145.06 241.16 ;
      RECT 144.8 240.92 149.4 241.08 ;
      RECT 135.8 240.92 143.38 241.08 ;
      RECT 135.8 239.96 149.4 240.12 ;
      RECT 135.8 242.4 149.4 242.56 ;
      RECT 144.8 241.36 145.06 242.56 ;
      RECT 144.8 241.44 149.4 241.6 ;
      RECT 135.8 241.44 143.38 241.6 ;
      RECT 143.1 241.36 145.06 241.52 ;
      RECT 143.1 244.4 145.06 244.56 ;
      RECT 144.8 243.36 145.06 244.56 ;
      RECT 144.8 244.32 149.4 244.48 ;
      RECT 135.8 244.32 143.38 244.48 ;
      RECT 135.8 243.36 149.4 243.52 ;
      RECT 135.8 245.8 149.4 245.96 ;
      RECT 144.8 244.76 145.06 245.96 ;
      RECT 144.8 244.84 149.4 245 ;
      RECT 135.8 244.84 143.38 245 ;
      RECT 143.1 244.76 145.06 244.92 ;
      RECT 143.1 247.8 145.06 247.96 ;
      RECT 144.8 246.76 145.06 247.96 ;
      RECT 144.8 247.72 149.4 247.88 ;
      RECT 135.8 247.72 143.38 247.88 ;
      RECT 135.8 246.76 149.4 246.92 ;
      RECT 135.8 249.2 149.4 249.36 ;
      RECT 144.8 248.16 145.06 249.36 ;
      RECT 144.8 248.24 149.4 248.4 ;
      RECT 135.8 248.24 143.38 248.4 ;
      RECT 143.1 248.16 145.06 248.32 ;
      RECT 143.1 251.2 145.06 251.36 ;
      RECT 144.8 250.16 145.06 251.36 ;
      RECT 144.8 251.12 149.4 251.28 ;
      RECT 135.8 251.12 143.38 251.28 ;
      RECT 135.8 250.16 149.4 250.32 ;
      RECT 135.8 252.6 149.4 252.76 ;
      RECT 144.8 251.56 145.06 252.76 ;
      RECT 144.8 251.64 149.4 251.8 ;
      RECT 135.8 251.64 143.38 251.8 ;
      RECT 143.1 251.56 145.06 251.72 ;
      RECT 143.1 254.6 145.06 254.76 ;
      RECT 144.8 253.56 145.06 254.76 ;
      RECT 144.8 254.52 149.4 254.68 ;
      RECT 135.8 254.52 143.38 254.68 ;
      RECT 135.8 253.56 149.4 253.72 ;
      RECT 135.8 256 149.4 256.16 ;
      RECT 144.8 254.96 145.06 256.16 ;
      RECT 144.8 255.04 149.4 255.2 ;
      RECT 135.8 255.04 143.38 255.2 ;
      RECT 143.1 254.96 145.06 255.12 ;
      RECT 143.1 258 145.06 258.16 ;
      RECT 144.8 256.96 145.06 258.16 ;
      RECT 144.8 257.92 149.4 258.08 ;
      RECT 135.8 257.92 143.38 258.08 ;
      RECT 135.8 256.96 149.4 257.12 ;
      RECT 135.8 259.4 149.4 259.56 ;
      RECT 144.8 258.36 145.06 259.56 ;
      RECT 144.8 258.44 149.4 258.6 ;
      RECT 135.8 258.44 143.38 258.6 ;
      RECT 143.1 258.36 145.06 258.52 ;
      RECT 143.1 261.4 145.06 261.56 ;
      RECT 144.8 260.36 145.06 261.56 ;
      RECT 144.8 261.32 149.4 261.48 ;
      RECT 135.8 261.32 143.38 261.48 ;
      RECT 135.8 260.36 149.4 260.52 ;
      RECT 135.8 262.8 149.4 262.96 ;
      RECT 144.8 261.76 145.06 262.96 ;
      RECT 144.8 261.84 149.4 262 ;
      RECT 135.8 261.84 143.38 262 ;
      RECT 143.1 261.76 145.06 261.92 ;
      RECT 143.1 264.8 145.06 264.96 ;
      RECT 144.8 263.76 145.06 264.96 ;
      RECT 144.8 264.72 149.4 264.88 ;
      RECT 135.8 264.72 143.38 264.88 ;
      RECT 135.8 263.76 149.4 263.92 ;
      RECT 135.8 266.2 149.4 266.36 ;
      RECT 144.8 265.16 145.06 266.36 ;
      RECT 144.8 265.24 149.4 265.4 ;
      RECT 135.8 265.24 143.38 265.4 ;
      RECT 143.1 265.16 145.06 265.32 ;
      RECT 143.1 268.2 145.06 268.36 ;
      RECT 144.8 267.16 145.06 268.36 ;
      RECT 144.8 268.12 149.4 268.28 ;
      RECT 135.8 268.12 143.38 268.28 ;
      RECT 135.8 267.16 149.4 267.32 ;
      RECT 135.8 269.6 149.4 269.76 ;
      RECT 144.8 268.56 145.06 269.76 ;
      RECT 144.8 268.64 149.4 268.8 ;
      RECT 135.8 268.64 143.38 268.8 ;
      RECT 143.1 268.56 145.06 268.72 ;
      RECT 143.1 271.6 145.06 271.76 ;
      RECT 144.8 270.56 145.06 271.76 ;
      RECT 144.8 271.52 149.4 271.68 ;
      RECT 135.8 271.52 143.38 271.68 ;
      RECT 135.8 270.56 149.4 270.72 ;
      RECT 135.8 273 149.4 273.16 ;
      RECT 144.8 271.96 145.06 273.16 ;
      RECT 144.8 272.04 149.4 272.2 ;
      RECT 135.8 272.04 143.38 272.2 ;
      RECT 143.1 271.96 145.06 272.12 ;
      RECT 143.1 275 145.06 275.16 ;
      RECT 144.8 273.96 145.06 275.16 ;
      RECT 144.8 274.92 149.4 275.08 ;
      RECT 135.8 274.92 143.38 275.08 ;
      RECT 135.8 273.96 149.4 274.12 ;
      RECT 135.8 276.4 149.4 276.56 ;
      RECT 144.8 275.36 145.06 276.56 ;
      RECT 144.8 275.44 149.4 275.6 ;
      RECT 135.8 275.44 143.38 275.6 ;
      RECT 143.1 275.36 145.06 275.52 ;
      RECT 143.1 278.4 145.06 278.56 ;
      RECT 144.8 277.36 145.06 278.56 ;
      RECT 144.8 278.32 149.4 278.48 ;
      RECT 135.8 278.32 143.38 278.48 ;
      RECT 135.8 277.36 149.4 277.52 ;
      RECT 135.8 279.8 149.4 279.96 ;
      RECT 144.8 278.76 145.06 279.96 ;
      RECT 144.8 278.84 149.4 279 ;
      RECT 135.8 278.84 143.38 279 ;
      RECT 143.1 278.76 145.06 278.92 ;
      RECT 143.1 281.8 145.06 281.96 ;
      RECT 144.8 280.76 145.06 281.96 ;
      RECT 144.8 281.72 149.4 281.88 ;
      RECT 135.8 281.72 143.38 281.88 ;
      RECT 135.8 280.76 149.4 280.92 ;
      RECT 135.8 283.2 149.4 283.36 ;
      RECT 144.8 282.16 145.06 283.36 ;
      RECT 144.8 282.24 149.4 282.4 ;
      RECT 135.8 282.24 143.38 282.4 ;
      RECT 143.1 282.16 145.06 282.32 ;
      RECT 143.1 285.2 145.06 285.36 ;
      RECT 144.8 284.16 145.06 285.36 ;
      RECT 144.8 285.12 149.4 285.28 ;
      RECT 135.8 285.12 143.38 285.28 ;
      RECT 135.8 284.16 149.4 284.32 ;
      RECT 135.8 286.6 149.4 286.76 ;
      RECT 144.8 285.56 145.06 286.76 ;
      RECT 144.8 285.64 149.4 285.8 ;
      RECT 135.8 285.64 143.38 285.8 ;
      RECT 143.1 285.56 145.06 285.72 ;
      RECT 143.1 288.6 145.06 288.76 ;
      RECT 144.8 287.56 145.06 288.76 ;
      RECT 144.8 288.52 149.4 288.68 ;
      RECT 135.8 288.52 143.38 288.68 ;
      RECT 135.8 287.56 149.4 287.72 ;
      RECT 135.8 290 149.4 290.16 ;
      RECT 144.8 288.96 145.06 290.16 ;
      RECT 144.8 289.04 149.4 289.2 ;
      RECT 135.8 289.04 143.38 289.2 ;
      RECT 143.1 288.96 145.06 289.12 ;
      RECT 143.1 292 145.06 292.16 ;
      RECT 144.8 290.96 145.06 292.16 ;
      RECT 144.8 291.92 149.4 292.08 ;
      RECT 135.8 291.92 143.38 292.08 ;
      RECT 135.8 290.96 149.4 291.12 ;
      RECT 135.8 293.4 149.4 293.56 ;
      RECT 144.8 292.36 145.06 293.56 ;
      RECT 144.8 292.44 149.4 292.6 ;
      RECT 135.8 292.44 143.38 292.6 ;
      RECT 143.1 292.36 145.06 292.52 ;
      RECT 143.1 295.4 145.06 295.56 ;
      RECT 144.8 294.36 145.06 295.56 ;
      RECT 144.8 295.32 149.4 295.48 ;
      RECT 135.8 295.32 143.38 295.48 ;
      RECT 135.8 294.36 149.4 294.52 ;
      RECT 135.8 296.8 149.4 296.96 ;
      RECT 144.8 295.76 145.06 296.96 ;
      RECT 144.8 295.84 149.4 296 ;
      RECT 135.8 295.84 143.38 296 ;
      RECT 143.1 295.76 145.06 295.92 ;
      RECT 143.1 298.8 145.06 298.96 ;
      RECT 144.8 297.76 145.06 298.96 ;
      RECT 144.8 298.72 149.4 298.88 ;
      RECT 135.8 298.72 143.38 298.88 ;
      RECT 135.8 297.76 149.4 297.92 ;
      RECT 135.8 300.2 149.4 300.36 ;
      RECT 144.8 299.16 145.06 300.36 ;
      RECT 144.8 299.24 149.4 299.4 ;
      RECT 135.8 299.24 143.38 299.4 ;
      RECT 143.1 299.16 145.06 299.32 ;
      RECT 143.1 302.2 145.06 302.36 ;
      RECT 144.8 301.16 145.06 302.36 ;
      RECT 144.8 302.12 149.4 302.28 ;
      RECT 135.8 302.12 143.38 302.28 ;
      RECT 135.8 301.16 149.4 301.32 ;
      RECT 135.8 303.6 149.4 303.76 ;
      RECT 144.8 302.56 145.06 303.76 ;
      RECT 144.8 302.64 149.4 302.8 ;
      RECT 135.8 302.64 143.38 302.8 ;
      RECT 143.1 302.56 145.06 302.72 ;
      RECT 143.1 305.6 145.06 305.76 ;
      RECT 144.8 304.56 145.06 305.76 ;
      RECT 144.8 305.52 149.4 305.68 ;
      RECT 135.8 305.52 143.38 305.68 ;
      RECT 135.8 304.56 149.4 304.72 ;
      RECT 135.8 307 149.4 307.16 ;
      RECT 144.8 305.96 145.06 307.16 ;
      RECT 144.8 306.04 149.4 306.2 ;
      RECT 135.8 306.04 143.38 306.2 ;
      RECT 143.1 305.96 145.06 306.12 ;
      RECT 143.1 309 145.06 309.16 ;
      RECT 144.8 307.96 145.06 309.16 ;
      RECT 144.8 308.92 149.4 309.08 ;
      RECT 135.8 308.92 143.38 309.08 ;
      RECT 135.8 307.96 149.4 308.12 ;
      RECT 135.8 310.4 149.4 310.56 ;
      RECT 144.8 309.36 145.06 310.56 ;
      RECT 144.8 309.44 149.4 309.6 ;
      RECT 135.8 309.44 143.38 309.6 ;
      RECT 143.1 309.36 145.06 309.52 ;
      RECT 143.1 312.4 145.06 312.56 ;
      RECT 144.8 311.36 145.06 312.56 ;
      RECT 144.8 312.32 149.4 312.48 ;
      RECT 135.8 312.32 143.38 312.48 ;
      RECT 135.8 311.36 149.4 311.52 ;
      RECT 135.8 313.8 149.4 313.96 ;
      RECT 144.8 312.76 145.06 313.96 ;
      RECT 144.8 312.84 149.4 313 ;
      RECT 135.8 312.84 143.38 313 ;
      RECT 143.1 312.76 145.06 312.92 ;
      RECT 143.1 315.8 145.06 315.96 ;
      RECT 144.8 314.76 145.06 315.96 ;
      RECT 144.8 315.72 149.4 315.88 ;
      RECT 135.8 315.72 143.38 315.88 ;
      RECT 135.8 314.76 149.4 314.92 ;
      RECT 135.8 317.2 149.4 317.36 ;
      RECT 144.8 316.16 145.06 317.36 ;
      RECT 144.8 316.24 149.4 316.4 ;
      RECT 135.8 316.24 143.38 316.4 ;
      RECT 143.1 316.16 145.06 316.32 ;
      RECT 143.1 319.2 145.06 319.36 ;
      RECT 144.8 318.16 145.06 319.36 ;
      RECT 144.8 319.12 149.4 319.28 ;
      RECT 135.8 319.12 143.38 319.28 ;
      RECT 135.8 318.16 149.4 318.32 ;
      RECT 135.8 320.6 149.4 320.76 ;
      RECT 144.8 319.56 145.06 320.76 ;
      RECT 144.8 319.64 149.4 319.8 ;
      RECT 135.8 319.64 143.38 319.8 ;
      RECT 143.1 319.56 145.06 319.72 ;
      RECT 143.1 322.6 145.06 322.76 ;
      RECT 144.8 321.56 145.06 322.76 ;
      RECT 144.8 322.52 149.4 322.68 ;
      RECT 135.8 322.52 143.38 322.68 ;
      RECT 135.8 321.56 149.4 321.72 ;
      RECT 135.8 324 149.4 324.16 ;
      RECT 144.8 322.96 145.06 324.16 ;
      RECT 144.8 323.04 149.4 323.2 ;
      RECT 135.8 323.04 143.38 323.2 ;
      RECT 143.1 322.96 145.06 323.12 ;
      RECT 143.1 326 145.06 326.16 ;
      RECT 144.8 324.96 145.06 326.16 ;
      RECT 144.8 325.92 149.4 326.08 ;
      RECT 135.8 325.92 143.38 326.08 ;
      RECT 135.8 324.96 149.4 325.12 ;
      RECT 135.8 327.4 149.4 327.56 ;
      RECT 144.8 326.36 145.06 327.56 ;
      RECT 144.8 326.44 149.4 326.6 ;
      RECT 135.8 326.44 143.38 326.6 ;
      RECT 143.1 326.36 145.06 326.52 ;
      RECT 143.1 329.4 145.06 329.56 ;
      RECT 144.8 328.36 145.06 329.56 ;
      RECT 144.8 329.32 149.4 329.48 ;
      RECT 135.8 329.32 143.38 329.48 ;
      RECT 135.8 328.36 149.4 328.52 ;
      RECT 135.8 330.8 149.4 330.96 ;
      RECT 144.8 329.76 145.06 330.96 ;
      RECT 144.8 329.84 149.4 330 ;
      RECT 135.8 329.84 143.38 330 ;
      RECT 143.1 329.76 145.06 329.92 ;
      RECT 143.1 332.8 145.06 332.96 ;
      RECT 144.8 331.76 145.06 332.96 ;
      RECT 144.8 332.72 149.4 332.88 ;
      RECT 135.8 332.72 143.38 332.88 ;
      RECT 135.8 331.76 149.4 331.92 ;
      RECT 135.8 334.2 149.4 334.36 ;
      RECT 144.8 333.16 145.06 334.36 ;
      RECT 144.8 333.24 149.4 333.4 ;
      RECT 135.8 333.24 143.38 333.4 ;
      RECT 143.1 333.16 145.06 333.32 ;
      RECT 143.1 336.2 145.06 336.36 ;
      RECT 144.8 335.16 145.06 336.36 ;
      RECT 144.8 336.12 149.4 336.28 ;
      RECT 135.8 336.12 143.38 336.28 ;
      RECT 135.8 335.16 149.4 335.32 ;
      RECT 135.8 337.6 149.4 337.76 ;
      RECT 144.8 336.56 145.06 337.76 ;
      RECT 144.8 336.64 149.4 336.8 ;
      RECT 135.8 336.64 143.38 336.8 ;
      RECT 143.1 336.56 145.06 336.72 ;
      RECT 143.1 339.6 145.06 339.76 ;
      RECT 144.8 338.56 145.06 339.76 ;
      RECT 144.8 339.52 149.4 339.68 ;
      RECT 135.8 339.52 143.38 339.68 ;
      RECT 135.8 338.56 149.4 338.72 ;
      RECT 135.8 341 149.4 341.16 ;
      RECT 144.8 339.96 145.06 341.16 ;
      RECT 144.8 340.04 149.4 340.2 ;
      RECT 135.8 340.04 143.38 340.2 ;
      RECT 143.1 339.96 145.06 340.12 ;
      RECT 143.1 343 145.06 343.16 ;
      RECT 144.8 341.96 145.06 343.16 ;
      RECT 144.8 342.92 149.4 343.08 ;
      RECT 135.8 342.92 143.38 343.08 ;
      RECT 135.8 341.96 149.4 342.12 ;
      RECT 135.8 344.4 149.4 344.56 ;
      RECT 144.8 343.36 145.06 344.56 ;
      RECT 144.8 343.44 149.4 343.6 ;
      RECT 135.8 343.44 143.38 343.6 ;
      RECT 143.1 343.36 145.06 343.52 ;
      RECT 143.1 346.4 145.06 346.56 ;
      RECT 144.8 345.36 145.06 346.56 ;
      RECT 144.8 346.32 149.4 346.48 ;
      RECT 135.8 346.32 143.38 346.48 ;
      RECT 135.8 345.36 149.4 345.52 ;
      RECT 135.8 347.8 149.4 347.96 ;
      RECT 144.8 346.76 145.06 347.96 ;
      RECT 144.8 346.84 149.4 347 ;
      RECT 135.8 346.84 143.38 347 ;
      RECT 143.1 346.76 145.06 346.92 ;
      RECT 143.1 349.8 145.06 349.96 ;
      RECT 144.8 348.76 145.06 349.96 ;
      RECT 144.8 349.72 149.4 349.88 ;
      RECT 135.8 349.72 143.38 349.88 ;
      RECT 135.8 348.76 149.4 348.92 ;
      RECT 135.8 351.2 149.4 351.36 ;
      RECT 144.8 350.16 145.06 351.36 ;
      RECT 144.8 350.24 149.4 350.4 ;
      RECT 135.8 350.24 143.38 350.4 ;
      RECT 143.1 350.16 145.06 350.32 ;
      RECT 143.1 353.2 145.06 353.36 ;
      RECT 144.8 352.16 145.06 353.36 ;
      RECT 144.8 353.12 149.4 353.28 ;
      RECT 135.8 353.12 143.38 353.28 ;
      RECT 135.8 352.16 149.4 352.32 ;
      RECT 135.8 354.6 149.4 354.76 ;
      RECT 144.8 353.56 145.06 354.76 ;
      RECT 144.8 353.64 149.4 353.8 ;
      RECT 135.8 353.64 143.38 353.8 ;
      RECT 143.1 353.56 145.06 353.72 ;
      RECT 143.1 356.6 145.06 356.76 ;
      RECT 144.8 355.56 145.06 356.76 ;
      RECT 144.8 356.52 149.4 356.68 ;
      RECT 135.8 356.52 143.38 356.68 ;
      RECT 135.8 355.56 149.4 355.72 ;
      RECT 135.8 358 149.4 358.16 ;
      RECT 144.8 356.96 145.06 358.16 ;
      RECT 144.8 357.04 149.4 357.2 ;
      RECT 135.8 357.04 143.38 357.2 ;
      RECT 143.1 356.96 145.06 357.12 ;
      RECT 143.1 360 145.06 360.16 ;
      RECT 144.8 358.96 145.06 360.16 ;
      RECT 144.8 359.92 149.4 360.08 ;
      RECT 135.8 359.92 143.38 360.08 ;
      RECT 135.8 358.96 149.4 359.12 ;
      RECT 135.8 361.4 149.4 361.56 ;
      RECT 144.8 360.36 145.06 361.56 ;
      RECT 144.8 360.44 149.4 360.6 ;
      RECT 135.8 360.44 143.38 360.6 ;
      RECT 143.1 360.36 145.06 360.52 ;
      RECT 143.1 363.4 145.06 363.56 ;
      RECT 144.8 362.36 145.06 363.56 ;
      RECT 144.8 363.32 149.4 363.48 ;
      RECT 135.8 363.32 143.38 363.48 ;
      RECT 135.8 362.36 149.4 362.52 ;
      RECT 135.8 364.8 149.4 364.96 ;
      RECT 144.8 363.76 145.06 364.96 ;
      RECT 144.8 363.84 149.4 364 ;
      RECT 135.8 363.84 143.38 364 ;
      RECT 143.1 363.76 145.06 363.92 ;
      RECT 143.1 366.8 145.06 366.96 ;
      RECT 144.8 365.76 145.06 366.96 ;
      RECT 144.8 366.72 149.4 366.88 ;
      RECT 135.8 366.72 143.38 366.88 ;
      RECT 135.8 365.76 149.4 365.92 ;
      RECT 135.8 368.2 149.4 368.36 ;
      RECT 144.8 367.16 145.06 368.36 ;
      RECT 144.8 367.24 149.4 367.4 ;
      RECT 135.8 367.24 143.38 367.4 ;
      RECT 143.1 367.16 145.06 367.32 ;
      RECT 143.1 370.2 145.06 370.36 ;
      RECT 144.8 369.16 145.06 370.36 ;
      RECT 144.8 370.12 149.4 370.28 ;
      RECT 135.8 370.12 143.38 370.28 ;
      RECT 135.8 369.16 149.4 369.32 ;
      RECT 135.8 371.6 149.4 371.76 ;
      RECT 144.8 370.56 145.06 371.76 ;
      RECT 144.8 370.64 149.4 370.8 ;
      RECT 135.8 370.64 143.38 370.8 ;
      RECT 143.1 370.56 145.06 370.72 ;
      RECT 143.1 373.6 145.06 373.76 ;
      RECT 144.8 372.56 145.06 373.76 ;
      RECT 144.8 373.52 149.4 373.68 ;
      RECT 135.8 373.52 143.38 373.68 ;
      RECT 135.8 372.56 149.4 372.72 ;
      RECT 135.8 375 149.4 375.16 ;
      RECT 144.8 373.96 145.06 375.16 ;
      RECT 144.8 374.04 149.4 374.2 ;
      RECT 135.8 374.04 143.38 374.2 ;
      RECT 143.1 373.96 145.06 374.12 ;
      RECT 143.1 377 145.06 377.16 ;
      RECT 144.8 375.96 145.06 377.16 ;
      RECT 144.8 376.92 149.4 377.08 ;
      RECT 135.8 376.92 143.38 377.08 ;
      RECT 135.8 375.96 149.4 376.12 ;
      RECT 135.8 378.4 149.4 378.56 ;
      RECT 144.8 377.36 145.06 378.56 ;
      RECT 144.8 377.44 149.4 377.6 ;
      RECT 135.8 377.44 143.38 377.6 ;
      RECT 143.1 377.36 145.06 377.52 ;
      RECT 143.1 380.4 145.06 380.56 ;
      RECT 144.8 379.36 145.06 380.56 ;
      RECT 144.8 380.32 149.4 380.48 ;
      RECT 135.8 380.32 143.38 380.48 ;
      RECT 135.8 379.36 149.4 379.52 ;
      RECT 135.8 381.8 149.4 381.96 ;
      RECT 144.8 380.76 145.06 381.96 ;
      RECT 144.8 380.84 149.4 381 ;
      RECT 135.8 380.84 143.38 381 ;
      RECT 143.1 380.76 145.06 380.92 ;
      RECT 143.1 383.8 145.06 383.96 ;
      RECT 144.8 382.76 145.06 383.96 ;
      RECT 144.8 383.72 149.4 383.88 ;
      RECT 135.8 383.72 143.38 383.88 ;
      RECT 135.8 382.76 149.4 382.92 ;
      RECT 135.8 385.2 149.4 385.36 ;
      RECT 144.8 384.16 145.06 385.36 ;
      RECT 144.8 384.24 149.4 384.4 ;
      RECT 135.8 384.24 143.38 384.4 ;
      RECT 143.1 384.16 145.06 384.32 ;
      RECT 143.1 387.2 145.06 387.36 ;
      RECT 144.8 386.16 145.06 387.36 ;
      RECT 144.8 387.12 149.4 387.28 ;
      RECT 135.8 387.12 143.38 387.28 ;
      RECT 135.8 386.16 149.4 386.32 ;
      RECT 135.8 388.6 149.4 388.76 ;
      RECT 144.8 387.56 145.06 388.76 ;
      RECT 144.8 387.64 149.4 387.8 ;
      RECT 135.8 387.64 143.38 387.8 ;
      RECT 143.1 387.56 145.06 387.72 ;
      RECT 143.1 390.6 145.06 390.76 ;
      RECT 144.8 389.56 145.06 390.76 ;
      RECT 144.8 390.52 149.4 390.68 ;
      RECT 135.8 390.52 143.38 390.68 ;
      RECT 135.8 389.56 149.4 389.72 ;
      RECT 135.8 392 149.4 392.16 ;
      RECT 144.8 390.96 145.06 392.16 ;
      RECT 144.8 391.04 149.4 391.2 ;
      RECT 135.8 391.04 143.38 391.2 ;
      RECT 143.1 390.96 145.06 391.12 ;
      RECT 143.1 394 145.06 394.16 ;
      RECT 144.8 392.96 145.06 394.16 ;
      RECT 144.8 393.92 149.4 394.08 ;
      RECT 135.8 393.92 143.38 394.08 ;
      RECT 135.8 392.96 149.4 393.12 ;
      RECT 135.8 395.4 149.4 395.56 ;
      RECT 144.8 394.36 145.06 395.56 ;
      RECT 144.8 394.44 149.4 394.6 ;
      RECT 135.8 394.44 143.38 394.6 ;
      RECT 143.1 394.36 145.06 394.52 ;
      RECT 143.1 397.4 145.06 397.56 ;
      RECT 144.8 396.36 145.06 397.56 ;
      RECT 144.8 397.32 149.4 397.48 ;
      RECT 135.8 397.32 143.38 397.48 ;
      RECT 135.8 396.36 149.4 396.52 ;
      RECT 135.8 398.8 149.4 398.96 ;
      RECT 144.8 397.76 145.06 398.96 ;
      RECT 144.8 397.84 149.4 398 ;
      RECT 135.8 397.84 143.38 398 ;
      RECT 143.1 397.76 145.06 397.92 ;
      RECT 143.1 400.8 145.06 400.96 ;
      RECT 144.8 399.76 145.06 400.96 ;
      RECT 144.8 400.72 149.4 400.88 ;
      RECT 135.8 400.72 143.38 400.88 ;
      RECT 135.8 399.76 149.4 399.92 ;
      RECT 135.8 402.2 149.4 402.36 ;
      RECT 144.8 401.16 145.06 402.36 ;
      RECT 144.8 401.24 149.4 401.4 ;
      RECT 135.8 401.24 143.38 401.4 ;
      RECT 143.1 401.16 145.06 401.32 ;
      RECT 143.1 404.2 145.06 404.36 ;
      RECT 144.8 403.16 145.06 404.36 ;
      RECT 144.8 404.12 149.4 404.28 ;
      RECT 135.8 404.12 143.38 404.28 ;
      RECT 135.8 403.16 149.4 403.32 ;
      RECT 135.8 405.6 149.4 405.76 ;
      RECT 144.8 404.56 145.06 405.76 ;
      RECT 144.8 404.64 149.4 404.8 ;
      RECT 135.8 404.64 143.38 404.8 ;
      RECT 143.1 404.56 145.06 404.72 ;
      RECT 143.1 407.6 145.06 407.76 ;
      RECT 144.8 406.56 145.06 407.76 ;
      RECT 144.8 407.52 149.4 407.68 ;
      RECT 135.8 407.52 143.38 407.68 ;
      RECT 135.8 406.56 149.4 406.72 ;
      RECT 135.8 409 149.4 409.16 ;
      RECT 144.8 407.96 145.06 409.16 ;
      RECT 144.8 408.04 149.4 408.2 ;
      RECT 135.8 408.04 143.38 408.2 ;
      RECT 143.1 407.96 145.06 408.12 ;
      RECT 143.1 411 145.06 411.16 ;
      RECT 144.8 409.96 145.06 411.16 ;
      RECT 144.8 410.92 149.4 411.08 ;
      RECT 135.8 410.92 143.38 411.08 ;
      RECT 135.8 409.96 149.4 410.12 ;
      RECT 135.8 412.4 149.4 412.56 ;
      RECT 144.8 411.36 145.06 412.56 ;
      RECT 144.8 411.44 149.4 411.6 ;
      RECT 135.8 411.44 143.38 411.6 ;
      RECT 143.1 411.36 145.06 411.52 ;
      RECT 143.1 414.4 145.06 414.56 ;
      RECT 144.8 413.36 145.06 414.56 ;
      RECT 144.8 414.32 149.4 414.48 ;
      RECT 135.8 414.32 143.38 414.48 ;
      RECT 135.8 413.36 149.4 413.52 ;
      RECT 135.8 415.8 149.4 415.96 ;
      RECT 144.8 414.76 145.06 415.96 ;
      RECT 144.8 414.84 149.4 415 ;
      RECT 135.8 414.84 143.38 415 ;
      RECT 143.1 414.76 145.06 414.92 ;
      RECT 143.1 417.8 145.06 417.96 ;
      RECT 144.8 416.76 145.06 417.96 ;
      RECT 144.8 417.72 149.4 417.88 ;
      RECT 135.8 417.72 143.38 417.88 ;
      RECT 135.8 416.76 149.4 416.92 ;
      RECT 135.8 419.2 149.4 419.36 ;
      RECT 144.8 418.16 145.06 419.36 ;
      RECT 144.8 418.24 149.4 418.4 ;
      RECT 135.8 418.24 143.38 418.4 ;
      RECT 143.1 418.16 145.06 418.32 ;
      RECT 143.1 421.2 145.06 421.36 ;
      RECT 144.8 420.16 145.06 421.36 ;
      RECT 144.8 421.12 149.4 421.28 ;
      RECT 135.8 421.12 143.38 421.28 ;
      RECT 135.8 420.16 149.4 420.32 ;
      RECT 135.8 422.6 149.4 422.76 ;
      RECT 144.8 421.56 145.06 422.76 ;
      RECT 144.8 421.64 149.4 421.8 ;
      RECT 135.8 421.64 143.38 421.8 ;
      RECT 143.1 421.56 145.06 421.72 ;
      RECT 143.1 424.6 145.06 424.76 ;
      RECT 144.8 423.56 145.06 424.76 ;
      RECT 144.8 424.52 149.4 424.68 ;
      RECT 135.8 424.52 143.38 424.68 ;
      RECT 135.8 423.56 149.4 423.72 ;
      RECT 135.8 426 149.4 426.16 ;
      RECT 144.8 424.96 145.06 426.16 ;
      RECT 144.8 425.04 149.4 425.2 ;
      RECT 135.8 425.04 143.38 425.2 ;
      RECT 143.1 424.96 145.06 425.12 ;
      RECT 143.1 428 145.06 428.16 ;
      RECT 144.8 426.96 145.06 428.16 ;
      RECT 144.8 427.92 149.4 428.08 ;
      RECT 135.8 427.92 143.38 428.08 ;
      RECT 135.8 426.96 149.4 427.12 ;
      RECT 135.8 429.4 149.4 429.56 ;
      RECT 144.8 428.36 145.06 429.56 ;
      RECT 144.8 428.44 149.4 428.6 ;
      RECT 135.8 428.44 143.38 428.6 ;
      RECT 143.1 428.36 145.06 428.52 ;
      RECT 143.1 431.4 145.06 431.56 ;
      RECT 144.8 430.36 145.06 431.56 ;
      RECT 144.8 431.32 149.4 431.48 ;
      RECT 135.8 431.32 143.38 431.48 ;
      RECT 135.8 430.36 149.4 430.52 ;
      RECT 135.8 432.8 149.4 432.96 ;
      RECT 144.8 431.76 145.06 432.96 ;
      RECT 144.8 431.84 149.4 432 ;
      RECT 135.8 431.84 143.38 432 ;
      RECT 143.1 431.76 145.06 431.92 ;
      RECT 143.1 434.8 145.06 434.96 ;
      RECT 144.8 433.76 145.06 434.96 ;
      RECT 144.8 434.72 149.4 434.88 ;
      RECT 135.8 434.72 143.38 434.88 ;
      RECT 135.8 433.76 149.4 433.92 ;
      RECT 135.8 436.2 149.4 436.36 ;
      RECT 144.8 435.16 145.06 436.36 ;
      RECT 144.8 435.24 149.4 435.4 ;
      RECT 135.8 435.24 143.38 435.4 ;
      RECT 143.1 435.16 145.06 435.32 ;
      RECT 143.1 438.2 145.06 438.36 ;
      RECT 144.8 437.16 145.06 438.36 ;
      RECT 144.8 438.12 149.4 438.28 ;
      RECT 135.8 438.12 143.38 438.28 ;
      RECT 135.8 437.16 149.4 437.32 ;
      RECT 135.8 439.6 149.4 439.76 ;
      RECT 144.8 438.56 145.06 439.76 ;
      RECT 144.8 438.64 149.4 438.8 ;
      RECT 135.8 438.64 143.38 438.8 ;
      RECT 143.1 438.56 145.06 438.72 ;
      RECT 143.1 441.6 145.06 441.76 ;
      RECT 144.8 440.56 145.06 441.76 ;
      RECT 144.8 441.52 149.4 441.68 ;
      RECT 135.8 441.52 143.38 441.68 ;
      RECT 135.8 440.56 149.4 440.72 ;
      RECT 135.8 443 149.4 443.16 ;
      RECT 144.8 441.96 145.06 443.16 ;
      RECT 144.8 442.04 149.4 442.2 ;
      RECT 135.8 442.04 143.38 442.2 ;
      RECT 143.1 441.96 145.06 442.12 ;
      RECT 143.1 445 145.06 445.16 ;
      RECT 144.8 443.96 145.06 445.16 ;
      RECT 144.8 444.92 149.4 445.08 ;
      RECT 135.8 444.92 143.38 445.08 ;
      RECT 135.8 443.96 149.4 444.12 ;
      RECT 135.8 446.4 149.4 446.56 ;
      RECT 144.8 445.36 145.06 446.56 ;
      RECT 144.8 445.44 149.4 445.6 ;
      RECT 135.8 445.44 143.38 445.6 ;
      RECT 143.1 445.36 145.06 445.52 ;
      RECT 143.1 448.4 145.06 448.56 ;
      RECT 144.8 447.36 145.06 448.56 ;
      RECT 144.8 448.32 149.4 448.48 ;
      RECT 135.8 448.32 143.38 448.48 ;
      RECT 135.8 447.36 149.4 447.52 ;
      RECT 135.8 449.8 149.4 449.96 ;
      RECT 144.8 448.76 145.06 449.96 ;
      RECT 144.8 448.84 149.4 449 ;
      RECT 135.8 448.84 143.38 449 ;
      RECT 143.1 448.76 145.06 448.92 ;
      RECT 143.1 451.8 145.06 451.96 ;
      RECT 144.8 450.76 145.06 451.96 ;
      RECT 144.8 451.72 149.4 451.88 ;
      RECT 135.8 451.72 143.38 451.88 ;
      RECT 135.8 450.76 149.4 450.92 ;
      RECT 135.8 453.2 149.4 453.36 ;
      RECT 144.8 452.16 145.06 453.36 ;
      RECT 144.8 452.24 149.4 452.4 ;
      RECT 135.8 452.24 143.38 452.4 ;
      RECT 143.1 452.16 145.06 452.32 ;
      RECT 143.1 455.2 145.06 455.36 ;
      RECT 144.8 454.16 145.06 455.36 ;
      RECT 144.8 455.12 149.4 455.28 ;
      RECT 135.8 455.12 143.38 455.28 ;
      RECT 135.8 454.16 149.4 454.32 ;
      RECT 135.8 456.6 149.4 456.76 ;
      RECT 144.8 455.56 145.06 456.76 ;
      RECT 144.8 455.64 149.4 455.8 ;
      RECT 135.8 455.64 143.38 455.8 ;
      RECT 143.1 455.56 145.06 455.72 ;
      RECT 143.1 458.6 145.06 458.76 ;
      RECT 144.8 457.56 145.06 458.76 ;
      RECT 144.8 458.52 149.4 458.68 ;
      RECT 135.8 458.52 143.38 458.68 ;
      RECT 135.8 457.56 149.4 457.72 ;
      RECT 135.8 460 149.4 460.16 ;
      RECT 144.8 458.96 145.06 460.16 ;
      RECT 144.8 459.04 149.4 459.2 ;
      RECT 135.8 459.04 143.38 459.2 ;
      RECT 143.1 458.96 145.06 459.12 ;
      RECT 143.1 462 145.06 462.16 ;
      RECT 144.8 460.96 145.06 462.16 ;
      RECT 144.8 461.92 149.4 462.08 ;
      RECT 135.8 461.92 143.38 462.08 ;
      RECT 135.8 460.96 149.4 461.12 ;
      RECT 135.8 463.4 149.4 463.56 ;
      RECT 144.8 462.36 145.06 463.56 ;
      RECT 144.8 462.44 149.4 462.6 ;
      RECT 135.8 462.44 143.38 462.6 ;
      RECT 143.1 462.36 145.06 462.52 ;
      RECT 143.1 465.4 145.06 465.56 ;
      RECT 144.8 464.36 145.06 465.56 ;
      RECT 144.8 465.32 149.4 465.48 ;
      RECT 135.8 465.32 143.38 465.48 ;
      RECT 135.8 464.36 149.4 464.52 ;
      RECT 135.8 466.8 149.4 466.96 ;
      RECT 144.8 465.76 145.06 466.96 ;
      RECT 144.8 465.84 149.4 466 ;
      RECT 135.8 465.84 143.38 466 ;
      RECT 143.1 465.76 145.06 465.92 ;
      RECT 143.1 468.8 145.06 468.96 ;
      RECT 144.8 467.76 145.06 468.96 ;
      RECT 144.8 468.72 149.4 468.88 ;
      RECT 135.8 468.72 143.38 468.88 ;
      RECT 135.8 467.76 149.4 467.92 ;
      RECT 135.8 470.2 149.4 470.36 ;
      RECT 144.8 469.16 145.06 470.36 ;
      RECT 144.8 469.24 149.4 469.4 ;
      RECT 135.8 469.24 143.38 469.4 ;
      RECT 143.1 469.16 145.06 469.32 ;
      RECT 143.1 472.2 145.06 472.36 ;
      RECT 144.8 471.16 145.06 472.36 ;
      RECT 144.8 472.12 149.4 472.28 ;
      RECT 135.8 472.12 143.38 472.28 ;
      RECT 135.8 471.16 149.4 471.32 ;
      RECT 135.8 473.6 149.4 473.76 ;
      RECT 144.8 472.56 145.06 473.76 ;
      RECT 144.8 472.64 149.4 472.8 ;
      RECT 135.8 472.64 143.38 472.8 ;
      RECT 143.1 472.56 145.06 472.72 ;
      RECT 143.1 475.6 145.06 475.76 ;
      RECT 144.8 474.56 145.06 475.76 ;
      RECT 144.8 475.52 149.4 475.68 ;
      RECT 135.8 475.52 143.38 475.68 ;
      RECT 135.8 474.56 149.4 474.72 ;
      RECT 135.8 477 149.4 477.16 ;
      RECT 144.8 475.96 145.06 477.16 ;
      RECT 144.8 476.04 149.4 476.2 ;
      RECT 135.8 476.04 143.38 476.2 ;
      RECT 143.1 475.96 145.06 476.12 ;
      RECT 143.1 479 145.06 479.16 ;
      RECT 144.8 477.96 145.06 479.16 ;
      RECT 144.8 478.92 149.4 479.08 ;
      RECT 135.8 478.92 143.38 479.08 ;
      RECT 135.8 477.96 149.4 478.12 ;
      RECT 135.8 480.4 149.4 480.56 ;
      RECT 144.8 479.36 145.06 480.56 ;
      RECT 144.8 479.44 149.4 479.6 ;
      RECT 135.8 479.44 143.38 479.6 ;
      RECT 143.1 479.36 145.06 479.52 ;
      RECT 143.1 482.4 145.06 482.56 ;
      RECT 144.8 481.36 145.06 482.56 ;
      RECT 144.8 482.32 149.4 482.48 ;
      RECT 135.8 482.32 143.38 482.48 ;
      RECT 135.8 481.36 149.4 481.52 ;
      RECT 135.8 483.8 149.4 483.96 ;
      RECT 144.8 482.76 145.06 483.96 ;
      RECT 144.8 482.84 149.4 483 ;
      RECT 135.8 482.84 143.38 483 ;
      RECT 143.1 482.76 145.06 482.92 ;
      RECT 143.1 485.8 145.06 485.96 ;
      RECT 144.8 484.76 145.06 485.96 ;
      RECT 144.8 485.72 149.4 485.88 ;
      RECT 135.8 485.72 143.38 485.88 ;
      RECT 135.8 484.76 149.4 484.92 ;
      RECT 135.8 487.2 149.4 487.36 ;
      RECT 144.8 486.16 145.06 487.36 ;
      RECT 144.8 486.24 149.4 486.4 ;
      RECT 135.8 486.24 143.38 486.4 ;
      RECT 143.1 486.16 145.06 486.32 ;
      RECT 143.1 489.2 145.06 489.36 ;
      RECT 144.8 488.16 145.06 489.36 ;
      RECT 144.8 489.12 149.4 489.28 ;
      RECT 135.8 489.12 143.38 489.28 ;
      RECT 135.8 488.16 149.4 488.32 ;
      RECT 135.8 490.6 149.4 490.76 ;
      RECT 144.8 489.56 145.06 490.76 ;
      RECT 144.8 489.64 149.4 489.8 ;
      RECT 135.8 489.64 143.38 489.8 ;
      RECT 143.1 489.56 145.06 489.72 ;
      RECT 143.1 492.6 145.06 492.76 ;
      RECT 144.8 491.56 145.06 492.76 ;
      RECT 144.8 492.52 149.4 492.68 ;
      RECT 135.8 492.52 143.38 492.68 ;
      RECT 135.8 491.56 149.4 491.72 ;
      RECT 135.8 494 149.4 494.16 ;
      RECT 144.8 492.96 145.06 494.16 ;
      RECT 144.8 493.04 149.4 493.2 ;
      RECT 135.8 493.04 143.38 493.2 ;
      RECT 143.1 492.96 145.06 493.12 ;
      RECT 143.1 496 145.06 496.16 ;
      RECT 144.8 494.96 145.06 496.16 ;
      RECT 144.8 495.92 149.4 496.08 ;
      RECT 135.8 495.92 143.38 496.08 ;
      RECT 135.8 494.96 149.4 495.12 ;
      RECT 135.8 497.4 149.4 497.56 ;
      RECT 144.8 496.36 145.06 497.56 ;
      RECT 144.8 496.44 149.4 496.6 ;
      RECT 135.8 496.44 143.38 496.6 ;
      RECT 143.1 496.36 145.06 496.52 ;
      RECT 143.1 499.4 145.06 499.56 ;
      RECT 144.8 498.36 145.06 499.56 ;
      RECT 144.8 499.32 149.4 499.48 ;
      RECT 135.8 499.32 143.38 499.48 ;
      RECT 135.8 498.36 149.4 498.52 ;
      RECT 135.8 500.8 149.4 500.96 ;
      RECT 144.8 499.76 145.06 500.96 ;
      RECT 144.8 499.84 149.4 500 ;
      RECT 135.8 499.84 143.38 500 ;
      RECT 143.1 499.76 145.06 499.92 ;
      RECT 143.1 502.8 145.06 502.96 ;
      RECT 144.8 501.76 145.06 502.96 ;
      RECT 144.8 502.72 149.4 502.88 ;
      RECT 135.8 502.72 143.38 502.88 ;
      RECT 135.8 501.76 149.4 501.92 ;
      RECT 135.8 504.2 149.4 504.36 ;
      RECT 144.8 503.16 145.06 504.36 ;
      RECT 144.8 503.24 149.4 503.4 ;
      RECT 135.8 503.24 143.38 503.4 ;
      RECT 143.1 503.16 145.06 503.32 ;
      RECT 135.83 506.16 149.4 506.32 ;
      RECT 144.83 506.12 149.4 506.32 ;
      RECT 143.54 505.16 143.7 506.32 ;
      RECT 144.83 505.16 144.99 506.32 ;
      RECT 136.13 505.16 149.4 505.32 ;
      RECT 149.09 42.85 149.39 43.09 ;
      RECT 148.81 42.85 149.39 43.03 ;
      RECT 148.9 16.37 149.06 17.39 ;
      RECT 148.08 16.37 149.36 16.53 ;
      RECT 149.2 15.91 149.36 16.53 ;
      RECT 148.73 509.04 148.89 509.54 ;
      RECT 147.97 509.04 148.13 509.54 ;
      RECT 146.99 509.04 147.15 509.54 ;
      RECT 146.99 509.04 149.29 509.2 ;
      RECT 149.13 507.6 149.29 509.2 ;
      RECT 147.48 507.6 147.64 509.2 ;
      RECT 148.73 507.6 149.29 507.76 ;
      RECT 146.99 507.6 148.13 507.76 ;
      RECT 147.97 507.26 148.13 507.76 ;
      RECT 148.73 507.26 148.89 507.76 ;
      RECT 146.99 507.26 147.15 507.76 ;
      RECT 147.45 21.29 147.61 21.9 ;
      RECT 146.07 17.55 146.23 21.9 ;
      RECT 147.49 17.87 147.65 21.45 ;
      RECT 147.03 17.55 147.19 21.31 ;
      RECT 145.11 17.55 145.27 21.27 ;
      RECT 148.65 18.36 148.81 21.21 ;
      RECT 148.28 18.36 148.81 18.52 ;
      RECT 148.28 17.11 148.44 18.52 ;
      RECT 147.03 17.87 148.44 18.03 ;
      RECT 145.11 17.55 147.19 17.71 ;
      RECT 146.56 16.37 146.72 17.71 ;
      RECT 145.6 16.36 145.76 17.71 ;
      RECT 147.76 15.91 147.92 17.35 ;
      RECT 147.76 16.77 148.74 16.93 ;
      RECT 147.45 32.66 148.59 32.82 ;
      RECT 148.43 30.63 148.59 32.82 ;
      RECT 147.45 30.04 147.61 32.82 ;
      RECT 147.39 30.04 147.61 32.58 ;
      RECT 147.95 42.85 148.25 43.09 ;
      RECT 147.95 42.85 148.53 43.03 ;
      RECT 148.32 15.59 148.48 16.19 ;
      RECT 146.69 15.59 148.48 15.75 ;
      RECT 146.69 14.98 146.85 15.75 ;
      RECT 146.69 14.98 147.01 15.14 ;
      RECT 147.93 27.43 148.25 27.77 ;
      RECT 147.93 27.43 148.43 27.63 ;
      RECT 147.19 37.35 148.27 37.51 ;
      RECT 148.11 35.68 148.27 37.51 ;
      RECT 147.15 35.68 147.31 36.68 ;
      RECT 147.05 35.68 148.37 35.84 ;
      RECT 148.21 34.58 148.37 35.84 ;
      RECT 147.05 34.58 147.21 35.84 ;
      RECT 148.11 34.58 148.37 34.86 ;
      RECT 147.05 34.58 147.31 34.86 ;
      RECT 147.63 42.53 147.79 46.23 ;
      RECT 147.15 42.53 148.27 42.69 ;
      RECT 148.11 37.99 148.27 42.69 ;
      RECT 147.15 37.99 147.31 42.69 ;
      RECT 147.15 43.34 147.31 47.95 ;
      RECT 147.15 46.47 148.27 46.63 ;
      RECT 148.11 43.34 148.27 46.63 ;
      RECT 147.37 51.95 148.05 52.11 ;
      RECT 147.63 51.6 147.79 52.11 ;
      RECT 147.63 47.16 147.79 51.33 ;
      RECT 145.71 47.16 145.87 51.33 ;
      RECT 145.71 48.4 147.79 48.59 ;
      RECT 146.67 47.14 146.83 48.59 ;
      RECT 147.17 42.85 147.47 43.09 ;
      RECT 146.89 42.85 147.47 43.03 ;
      RECT 145.53 26.81 145.69 29.44 ;
      RECT 147.13 26.81 147.29 29.37 ;
      RECT 141.99 26.81 147.29 26.97 ;
      RECT 141.99 23.43 142.15 26.97 ;
      RECT 146.01 32.6 147.13 32.76 ;
      RECT 146.97 30.63 147.13 32.76 ;
      RECT 146.01 29.36 146.17 32.76 ;
      RECT 146.01 29.36 146.49 29.52 ;
      RECT 146.33 27.34 146.49 29.52 ;
      RECT 146.03 42.85 146.33 43.09 ;
      RECT 146.03 42.85 146.61 43.03 ;
      RECT 145.07 52.33 146.51 52.55 ;
      RECT 146.29 51.48 146.51 52.55 ;
      RECT 143.15 52.33 144.59 52.55 ;
      RECT 144.37 51.44 144.59 52.55 ;
      RECT 145.07 51.44 145.29 52.55 ;
      RECT 143.15 51.48 143.37 52.55 ;
      RECT 146.19 48.78 146.35 51.77 ;
      RECT 145.23 46.79 145.39 51.77 ;
      RECT 144.27 46.79 144.43 51.77 ;
      RECT 143.31 48.78 143.47 51.77 ;
      RECT 145.23 46.79 146.03 47 ;
      RECT 143.63 46.79 144.43 47 ;
      RECT 143.63 46.79 146.03 46.96 ;
      RECT 144.75 43.19 144.91 46.96 ;
      RECT 145.23 37.35 146.31 37.51 ;
      RECT 145.23 35.68 145.39 37.51 ;
      RECT 146.19 35.68 146.35 36.68 ;
      RECT 145.13 35.68 146.45 35.84 ;
      RECT 146.29 34.58 146.45 35.84 ;
      RECT 145.13 34.58 145.29 35.84 ;
      RECT 146.19 34.58 146.45 34.86 ;
      RECT 145.13 34.58 145.39 34.86 ;
      RECT 146.23 509.04 146.39 509.54 ;
      RECT 145.25 509.04 145.41 509.54 ;
      RECT 145.25 509.04 146.39 509.2 ;
      RECT 145.74 507.6 145.9 509.2 ;
      RECT 145.25 507.6 146.39 507.76 ;
      RECT 146.23 507.26 146.39 507.76 ;
      RECT 145.25 507.26 145.41 507.76 ;
      RECT 145.71 42.53 145.87 46.23 ;
      RECT 145.23 42.53 146.35 42.69 ;
      RECT 146.19 37.99 146.35 42.69 ;
      RECT 145.23 37.99 145.39 42.69 ;
      RECT 146.19 43.34 146.35 47.95 ;
      RECT 145.23 46.47 146.35 46.63 ;
      RECT 145.23 43.34 145.39 46.63 ;
      RECT 145.45 51.95 146.13 52.11 ;
      RECT 145.71 51.6 145.87 52.11 ;
      RECT 143.34 32.51 145.17 32.67 ;
      RECT 145.01 30.03 145.17 32.67 ;
      RECT 143.34 31.43 143.5 32.67 ;
      RECT 145.69 29.79 145.85 30.47 ;
      RECT 145.01 30.03 145.85 30.2 ;
      RECT 145.1 29.28 145.37 30.2 ;
      RECT 144.73 29.28 145.37 29.44 ;
      RECT 144.73 27.77 144.89 29.44 ;
      RECT 143.07 27.77 144.89 27.93 ;
      RECT 144.65 15.08 144.81 15.92 ;
      RECT 145.6 14.87 145.76 15.63 ;
      RECT 144.65 15.08 145.76 15.24 ;
      RECT 145.14 14.87 145.76 15.24 ;
      RECT 145.09 14.88 145.76 15.24 ;
      RECT 145.14 14.45 145.3 15.24 ;
      RECT 145.25 42.85 145.55 43.09 ;
      RECT 144.97 42.85 145.55 43.03 ;
      RECT 142.47 25.58 143.37 25.74 ;
      RECT 142.47 23.01 142.63 25.74 ;
      RECT 142.47 23.01 143.66 23.17 ;
      RECT 143.5 22.06 143.66 23.17 ;
      RECT 144.44 22.98 145.43 23.15 ;
      RECT 144.82 22.88 145.43 23.15 ;
      RECT 144.82 22.06 144.98 23.15 ;
      RECT 143.5 22.06 145.43 22.22 ;
      RECT 145.27 21.43 145.43 22.22 ;
      RECT 144.19 19.22 144.35 22.22 ;
      RECT 143.21 21.23 144.35 21.39 ;
      RECT 144.17 19.22 144.35 21.39 ;
      RECT 143.21 19.22 143.37 21.39 ;
      RECT 142.95 23.33 143.11 25.4 ;
      RECT 144.71 23.33 144.87 25.37 ;
      RECT 142.95 23.33 144.87 23.49 ;
      RECT 144.02 22.82 144.18 23.49 ;
      RECT 144.69 21.25 144.85 21.9 ;
      RECT 144.65 16.86 144.81 21.39 ;
      RECT 143.69 18.69 143.85 21.07 ;
      RECT 142.73 18.69 142.89 21.07 ;
      RECT 142.27 19.09 142.43 19.6 ;
      RECT 142.27 19.09 142.89 19.25 ;
      RECT 142.73 18.69 144.81 18.85 ;
      RECT 143.34 18.17 143.5 18.85 ;
      RECT 144.11 42.85 144.41 43.09 ;
      RECT 144.11 42.85 144.69 43.03 ;
      RECT 144.49 509.04 144.65 509.54 ;
      RECT 143.51 509.04 143.67 509.54 ;
      RECT 143.51 509.04 144.65 509.2 ;
      RECT 144 507.6 144.16 509.2 ;
      RECT 143.51 507.6 144.65 507.76 ;
      RECT 144.49 507.26 144.65 507.76 ;
      RECT 143.51 507.26 143.67 507.76 ;
      RECT 143.54 70.68 144.64 70.84 ;
      RECT 143.54 70.28 143.7 70.84 ;
      RECT 143.54 70.28 144.64 70.44 ;
      RECT 143.54 72.08 144.64 72.24 ;
      RECT 143.54 71.68 143.7 72.24 ;
      RECT 143.54 71.68 144.64 71.84 ;
      RECT 143.54 74.08 144.64 74.24 ;
      RECT 143.54 73.68 143.7 74.24 ;
      RECT 143.54 73.68 144.64 73.84 ;
      RECT 143.54 75.48 144.64 75.64 ;
      RECT 143.54 75.08 143.7 75.64 ;
      RECT 143.54 75.08 144.64 75.24 ;
      RECT 143.54 77.48 144.64 77.64 ;
      RECT 143.54 77.08 143.7 77.64 ;
      RECT 143.54 77.08 144.64 77.24 ;
      RECT 143.54 78.88 144.64 79.04 ;
      RECT 143.54 78.48 143.7 79.04 ;
      RECT 143.54 78.48 144.64 78.64 ;
      RECT 143.54 80.88 144.64 81.04 ;
      RECT 143.54 80.48 143.7 81.04 ;
      RECT 143.54 80.48 144.64 80.64 ;
      RECT 143.54 82.28 144.64 82.44 ;
      RECT 143.54 81.88 143.7 82.44 ;
      RECT 143.54 81.88 144.64 82.04 ;
      RECT 143.54 84.28 144.64 84.44 ;
      RECT 143.54 83.88 143.7 84.44 ;
      RECT 143.54 83.88 144.64 84.04 ;
      RECT 143.54 85.68 144.64 85.84 ;
      RECT 143.54 85.28 143.7 85.84 ;
      RECT 143.54 85.28 144.64 85.44 ;
      RECT 143.54 87.68 144.64 87.84 ;
      RECT 143.54 87.28 143.7 87.84 ;
      RECT 143.54 87.28 144.64 87.44 ;
      RECT 143.54 89.08 144.64 89.24 ;
      RECT 143.54 88.68 143.7 89.24 ;
      RECT 143.54 88.68 144.64 88.84 ;
      RECT 143.54 91.08 144.64 91.24 ;
      RECT 143.54 90.68 143.7 91.24 ;
      RECT 143.54 90.68 144.64 90.84 ;
      RECT 143.54 92.48 144.64 92.64 ;
      RECT 143.54 92.08 143.7 92.64 ;
      RECT 143.54 92.08 144.64 92.24 ;
      RECT 143.54 94.48 144.64 94.64 ;
      RECT 143.54 94.08 143.7 94.64 ;
      RECT 143.54 94.08 144.64 94.24 ;
      RECT 143.54 95.88 144.64 96.04 ;
      RECT 143.54 95.48 143.7 96.04 ;
      RECT 143.54 95.48 144.64 95.64 ;
      RECT 143.54 97.88 144.64 98.04 ;
      RECT 143.54 97.48 143.7 98.04 ;
      RECT 143.54 97.48 144.64 97.64 ;
      RECT 143.54 99.28 144.64 99.44 ;
      RECT 143.54 98.88 143.7 99.44 ;
      RECT 143.54 98.88 144.64 99.04 ;
      RECT 143.54 101.28 144.64 101.44 ;
      RECT 143.54 100.88 143.7 101.44 ;
      RECT 143.54 100.88 144.64 101.04 ;
      RECT 143.54 102.68 144.64 102.84 ;
      RECT 143.54 102.28 143.7 102.84 ;
      RECT 143.54 102.28 144.64 102.44 ;
      RECT 143.54 104.68 144.64 104.84 ;
      RECT 143.54 104.28 143.7 104.84 ;
      RECT 143.54 104.28 144.64 104.44 ;
      RECT 143.54 106.08 144.64 106.24 ;
      RECT 143.54 105.68 143.7 106.24 ;
      RECT 143.54 105.68 144.64 105.84 ;
      RECT 143.54 108.08 144.64 108.24 ;
      RECT 143.54 107.68 143.7 108.24 ;
      RECT 143.54 107.68 144.64 107.84 ;
      RECT 143.54 109.48 144.64 109.64 ;
      RECT 143.54 109.08 143.7 109.64 ;
      RECT 143.54 109.08 144.64 109.24 ;
      RECT 143.54 111.48 144.64 111.64 ;
      RECT 143.54 111.08 143.7 111.64 ;
      RECT 143.54 111.08 144.64 111.24 ;
      RECT 143.54 112.88 144.64 113.04 ;
      RECT 143.54 112.48 143.7 113.04 ;
      RECT 143.54 112.48 144.64 112.64 ;
      RECT 143.54 114.88 144.64 115.04 ;
      RECT 143.54 114.48 143.7 115.04 ;
      RECT 143.54 114.48 144.64 114.64 ;
      RECT 143.54 116.28 144.64 116.44 ;
      RECT 143.54 115.88 143.7 116.44 ;
      RECT 143.54 115.88 144.64 116.04 ;
      RECT 143.54 118.28 144.64 118.44 ;
      RECT 143.54 117.88 143.7 118.44 ;
      RECT 143.54 117.88 144.64 118.04 ;
      RECT 143.54 119.68 144.64 119.84 ;
      RECT 143.54 119.28 143.7 119.84 ;
      RECT 143.54 119.28 144.64 119.44 ;
      RECT 143.54 121.68 144.64 121.84 ;
      RECT 143.54 121.28 143.7 121.84 ;
      RECT 143.54 121.28 144.64 121.44 ;
      RECT 143.54 123.08 144.64 123.24 ;
      RECT 143.54 122.68 143.7 123.24 ;
      RECT 143.54 122.68 144.64 122.84 ;
      RECT 143.54 125.08 144.64 125.24 ;
      RECT 143.54 124.68 143.7 125.24 ;
      RECT 143.54 124.68 144.64 124.84 ;
      RECT 143.54 126.48 144.64 126.64 ;
      RECT 143.54 126.08 143.7 126.64 ;
      RECT 143.54 126.08 144.64 126.24 ;
      RECT 143.54 128.48 144.64 128.64 ;
      RECT 143.54 128.08 143.7 128.64 ;
      RECT 143.54 128.08 144.64 128.24 ;
      RECT 143.54 129.88 144.64 130.04 ;
      RECT 143.54 129.48 143.7 130.04 ;
      RECT 143.54 129.48 144.64 129.64 ;
      RECT 143.54 131.88 144.64 132.04 ;
      RECT 143.54 131.48 143.7 132.04 ;
      RECT 143.54 131.48 144.64 131.64 ;
      RECT 143.54 133.28 144.64 133.44 ;
      RECT 143.54 132.88 143.7 133.44 ;
      RECT 143.54 132.88 144.64 133.04 ;
      RECT 143.54 135.28 144.64 135.44 ;
      RECT 143.54 134.88 143.7 135.44 ;
      RECT 143.54 134.88 144.64 135.04 ;
      RECT 143.54 136.68 144.64 136.84 ;
      RECT 143.54 136.28 143.7 136.84 ;
      RECT 143.54 136.28 144.64 136.44 ;
      RECT 143.54 138.68 144.64 138.84 ;
      RECT 143.54 138.28 143.7 138.84 ;
      RECT 143.54 138.28 144.64 138.44 ;
      RECT 143.54 140.08 144.64 140.24 ;
      RECT 143.54 139.68 143.7 140.24 ;
      RECT 143.54 139.68 144.64 139.84 ;
      RECT 143.54 142.08 144.64 142.24 ;
      RECT 143.54 141.68 143.7 142.24 ;
      RECT 143.54 141.68 144.64 141.84 ;
      RECT 143.54 143.48 144.64 143.64 ;
      RECT 143.54 143.08 143.7 143.64 ;
      RECT 143.54 143.08 144.64 143.24 ;
      RECT 143.54 145.48 144.64 145.64 ;
      RECT 143.54 145.08 143.7 145.64 ;
      RECT 143.54 145.08 144.64 145.24 ;
      RECT 143.54 146.88 144.64 147.04 ;
      RECT 143.54 146.48 143.7 147.04 ;
      RECT 143.54 146.48 144.64 146.64 ;
      RECT 143.54 148.88 144.64 149.04 ;
      RECT 143.54 148.48 143.7 149.04 ;
      RECT 143.54 148.48 144.64 148.64 ;
      RECT 143.54 150.28 144.64 150.44 ;
      RECT 143.54 149.88 143.7 150.44 ;
      RECT 143.54 149.88 144.64 150.04 ;
      RECT 143.54 152.28 144.64 152.44 ;
      RECT 143.54 151.88 143.7 152.44 ;
      RECT 143.54 151.88 144.64 152.04 ;
      RECT 143.54 153.68 144.64 153.84 ;
      RECT 143.54 153.28 143.7 153.84 ;
      RECT 143.54 153.28 144.64 153.44 ;
      RECT 143.54 155.68 144.64 155.84 ;
      RECT 143.54 155.28 143.7 155.84 ;
      RECT 143.54 155.28 144.64 155.44 ;
      RECT 143.54 157.08 144.64 157.24 ;
      RECT 143.54 156.68 143.7 157.24 ;
      RECT 143.54 156.68 144.64 156.84 ;
      RECT 143.54 159.08 144.64 159.24 ;
      RECT 143.54 158.68 143.7 159.24 ;
      RECT 143.54 158.68 144.64 158.84 ;
      RECT 143.54 160.48 144.64 160.64 ;
      RECT 143.54 160.08 143.7 160.64 ;
      RECT 143.54 160.08 144.64 160.24 ;
      RECT 143.54 162.48 144.64 162.64 ;
      RECT 143.54 162.08 143.7 162.64 ;
      RECT 143.54 162.08 144.64 162.24 ;
      RECT 143.54 163.88 144.64 164.04 ;
      RECT 143.54 163.48 143.7 164.04 ;
      RECT 143.54 163.48 144.64 163.64 ;
      RECT 143.54 165.88 144.64 166.04 ;
      RECT 143.54 165.48 143.7 166.04 ;
      RECT 143.54 165.48 144.64 165.64 ;
      RECT 143.54 167.28 144.64 167.44 ;
      RECT 143.54 166.88 143.7 167.44 ;
      RECT 143.54 166.88 144.64 167.04 ;
      RECT 143.54 169.28 144.64 169.44 ;
      RECT 143.54 168.88 143.7 169.44 ;
      RECT 143.54 168.88 144.64 169.04 ;
      RECT 143.54 170.68 144.64 170.84 ;
      RECT 143.54 170.28 143.7 170.84 ;
      RECT 143.54 170.28 144.64 170.44 ;
      RECT 143.54 172.68 144.64 172.84 ;
      RECT 143.54 172.28 143.7 172.84 ;
      RECT 143.54 172.28 144.64 172.44 ;
      RECT 143.54 174.08 144.64 174.24 ;
      RECT 143.54 173.68 143.7 174.24 ;
      RECT 143.54 173.68 144.64 173.84 ;
      RECT 143.54 176.08 144.64 176.24 ;
      RECT 143.54 175.68 143.7 176.24 ;
      RECT 143.54 175.68 144.64 175.84 ;
      RECT 143.54 177.48 144.64 177.64 ;
      RECT 143.54 177.08 143.7 177.64 ;
      RECT 143.54 177.08 144.64 177.24 ;
      RECT 143.54 179.48 144.64 179.64 ;
      RECT 143.54 179.08 143.7 179.64 ;
      RECT 143.54 179.08 144.64 179.24 ;
      RECT 143.54 180.88 144.64 181.04 ;
      RECT 143.54 180.48 143.7 181.04 ;
      RECT 143.54 180.48 144.64 180.64 ;
      RECT 143.54 182.88 144.64 183.04 ;
      RECT 143.54 182.48 143.7 183.04 ;
      RECT 143.54 182.48 144.64 182.64 ;
      RECT 143.54 184.28 144.64 184.44 ;
      RECT 143.54 183.88 143.7 184.44 ;
      RECT 143.54 183.88 144.64 184.04 ;
      RECT 143.54 186.28 144.64 186.44 ;
      RECT 143.54 185.88 143.7 186.44 ;
      RECT 143.54 185.88 144.64 186.04 ;
      RECT 143.54 187.68 144.64 187.84 ;
      RECT 143.54 187.28 143.7 187.84 ;
      RECT 143.54 187.28 144.64 187.44 ;
      RECT 143.54 189.68 144.64 189.84 ;
      RECT 143.54 189.28 143.7 189.84 ;
      RECT 143.54 189.28 144.64 189.44 ;
      RECT 143.54 191.08 144.64 191.24 ;
      RECT 143.54 190.68 143.7 191.24 ;
      RECT 143.54 190.68 144.64 190.84 ;
      RECT 143.54 193.08 144.64 193.24 ;
      RECT 143.54 192.68 143.7 193.24 ;
      RECT 143.54 192.68 144.64 192.84 ;
      RECT 143.54 194.48 144.64 194.64 ;
      RECT 143.54 194.08 143.7 194.64 ;
      RECT 143.54 194.08 144.64 194.24 ;
      RECT 143.54 196.48 144.64 196.64 ;
      RECT 143.54 196.08 143.7 196.64 ;
      RECT 143.54 196.08 144.64 196.24 ;
      RECT 143.54 197.88 144.64 198.04 ;
      RECT 143.54 197.48 143.7 198.04 ;
      RECT 143.54 197.48 144.64 197.64 ;
      RECT 143.54 199.88 144.64 200.04 ;
      RECT 143.54 199.48 143.7 200.04 ;
      RECT 143.54 199.48 144.64 199.64 ;
      RECT 143.54 201.28 144.64 201.44 ;
      RECT 143.54 200.88 143.7 201.44 ;
      RECT 143.54 200.88 144.64 201.04 ;
      RECT 143.54 203.28 144.64 203.44 ;
      RECT 143.54 202.88 143.7 203.44 ;
      RECT 143.54 202.88 144.64 203.04 ;
      RECT 143.54 204.68 144.64 204.84 ;
      RECT 143.54 204.28 143.7 204.84 ;
      RECT 143.54 204.28 144.64 204.44 ;
      RECT 143.54 206.68 144.64 206.84 ;
      RECT 143.54 206.28 143.7 206.84 ;
      RECT 143.54 206.28 144.64 206.44 ;
      RECT 143.54 208.08 144.64 208.24 ;
      RECT 143.54 207.68 143.7 208.24 ;
      RECT 143.54 207.68 144.64 207.84 ;
      RECT 143.54 210.08 144.64 210.24 ;
      RECT 143.54 209.68 143.7 210.24 ;
      RECT 143.54 209.68 144.64 209.84 ;
      RECT 143.54 211.48 144.64 211.64 ;
      RECT 143.54 211.08 143.7 211.64 ;
      RECT 143.54 211.08 144.64 211.24 ;
      RECT 143.54 213.48 144.64 213.64 ;
      RECT 143.54 213.08 143.7 213.64 ;
      RECT 143.54 213.08 144.64 213.24 ;
      RECT 143.54 214.88 144.64 215.04 ;
      RECT 143.54 214.48 143.7 215.04 ;
      RECT 143.54 214.48 144.64 214.64 ;
      RECT 143.54 216.88 144.64 217.04 ;
      RECT 143.54 216.48 143.7 217.04 ;
      RECT 143.54 216.48 144.64 216.64 ;
      RECT 143.54 218.28 144.64 218.44 ;
      RECT 143.54 217.88 143.7 218.44 ;
      RECT 143.54 217.88 144.64 218.04 ;
      RECT 143.54 220.28 144.64 220.44 ;
      RECT 143.54 219.88 143.7 220.44 ;
      RECT 143.54 219.88 144.64 220.04 ;
      RECT 143.54 221.68 144.64 221.84 ;
      RECT 143.54 221.28 143.7 221.84 ;
      RECT 143.54 221.28 144.64 221.44 ;
      RECT 143.54 223.68 144.64 223.84 ;
      RECT 143.54 223.28 143.7 223.84 ;
      RECT 143.54 223.28 144.64 223.44 ;
      RECT 143.54 225.08 144.64 225.24 ;
      RECT 143.54 224.68 143.7 225.24 ;
      RECT 143.54 224.68 144.64 224.84 ;
      RECT 143.54 227.08 144.64 227.24 ;
      RECT 143.54 226.68 143.7 227.24 ;
      RECT 143.54 226.68 144.64 226.84 ;
      RECT 143.54 228.48 144.64 228.64 ;
      RECT 143.54 228.08 143.7 228.64 ;
      RECT 143.54 228.08 144.64 228.24 ;
      RECT 143.54 230.48 144.64 230.64 ;
      RECT 143.54 230.08 143.7 230.64 ;
      RECT 143.54 230.08 144.64 230.24 ;
      RECT 143.54 231.88 144.64 232.04 ;
      RECT 143.54 231.48 143.7 232.04 ;
      RECT 143.54 231.48 144.64 231.64 ;
      RECT 143.54 233.88 144.64 234.04 ;
      RECT 143.54 233.48 143.7 234.04 ;
      RECT 143.54 233.48 144.64 233.64 ;
      RECT 143.54 235.28 144.64 235.44 ;
      RECT 143.54 234.88 143.7 235.44 ;
      RECT 143.54 234.88 144.64 235.04 ;
      RECT 143.54 237.28 144.64 237.44 ;
      RECT 143.54 236.88 143.7 237.44 ;
      RECT 143.54 236.88 144.64 237.04 ;
      RECT 143.54 238.68 144.64 238.84 ;
      RECT 143.54 238.28 143.7 238.84 ;
      RECT 143.54 238.28 144.64 238.44 ;
      RECT 143.54 240.68 144.64 240.84 ;
      RECT 143.54 240.28 143.7 240.84 ;
      RECT 143.54 240.28 144.64 240.44 ;
      RECT 143.54 242.08 144.64 242.24 ;
      RECT 143.54 241.68 143.7 242.24 ;
      RECT 143.54 241.68 144.64 241.84 ;
      RECT 143.54 244.08 144.64 244.24 ;
      RECT 143.54 243.68 143.7 244.24 ;
      RECT 143.54 243.68 144.64 243.84 ;
      RECT 143.54 245.48 144.64 245.64 ;
      RECT 143.54 245.08 143.7 245.64 ;
      RECT 143.54 245.08 144.64 245.24 ;
      RECT 143.54 247.48 144.64 247.64 ;
      RECT 143.54 247.08 143.7 247.64 ;
      RECT 143.54 247.08 144.64 247.24 ;
      RECT 143.54 248.88 144.64 249.04 ;
      RECT 143.54 248.48 143.7 249.04 ;
      RECT 143.54 248.48 144.64 248.64 ;
      RECT 143.54 250.88 144.64 251.04 ;
      RECT 143.54 250.48 143.7 251.04 ;
      RECT 143.54 250.48 144.64 250.64 ;
      RECT 143.54 252.28 144.64 252.44 ;
      RECT 143.54 251.88 143.7 252.44 ;
      RECT 143.54 251.88 144.64 252.04 ;
      RECT 143.54 254.28 144.64 254.44 ;
      RECT 143.54 253.88 143.7 254.44 ;
      RECT 143.54 253.88 144.64 254.04 ;
      RECT 143.54 255.68 144.64 255.84 ;
      RECT 143.54 255.28 143.7 255.84 ;
      RECT 143.54 255.28 144.64 255.44 ;
      RECT 143.54 257.68 144.64 257.84 ;
      RECT 143.54 257.28 143.7 257.84 ;
      RECT 143.54 257.28 144.64 257.44 ;
      RECT 143.54 259.08 144.64 259.24 ;
      RECT 143.54 258.68 143.7 259.24 ;
      RECT 143.54 258.68 144.64 258.84 ;
      RECT 143.54 261.08 144.64 261.24 ;
      RECT 143.54 260.68 143.7 261.24 ;
      RECT 143.54 260.68 144.64 260.84 ;
      RECT 143.54 262.48 144.64 262.64 ;
      RECT 143.54 262.08 143.7 262.64 ;
      RECT 143.54 262.08 144.64 262.24 ;
      RECT 143.54 264.48 144.64 264.64 ;
      RECT 143.54 264.08 143.7 264.64 ;
      RECT 143.54 264.08 144.64 264.24 ;
      RECT 143.54 265.88 144.64 266.04 ;
      RECT 143.54 265.48 143.7 266.04 ;
      RECT 143.54 265.48 144.64 265.64 ;
      RECT 143.54 267.88 144.64 268.04 ;
      RECT 143.54 267.48 143.7 268.04 ;
      RECT 143.54 267.48 144.64 267.64 ;
      RECT 143.54 269.28 144.64 269.44 ;
      RECT 143.54 268.88 143.7 269.44 ;
      RECT 143.54 268.88 144.64 269.04 ;
      RECT 143.54 271.28 144.64 271.44 ;
      RECT 143.54 270.88 143.7 271.44 ;
      RECT 143.54 270.88 144.64 271.04 ;
      RECT 143.54 272.68 144.64 272.84 ;
      RECT 143.54 272.28 143.7 272.84 ;
      RECT 143.54 272.28 144.64 272.44 ;
      RECT 143.54 274.68 144.64 274.84 ;
      RECT 143.54 274.28 143.7 274.84 ;
      RECT 143.54 274.28 144.64 274.44 ;
      RECT 143.54 276.08 144.64 276.24 ;
      RECT 143.54 275.68 143.7 276.24 ;
      RECT 143.54 275.68 144.64 275.84 ;
      RECT 143.54 278.08 144.64 278.24 ;
      RECT 143.54 277.68 143.7 278.24 ;
      RECT 143.54 277.68 144.64 277.84 ;
      RECT 143.54 279.48 144.64 279.64 ;
      RECT 143.54 279.08 143.7 279.64 ;
      RECT 143.54 279.08 144.64 279.24 ;
      RECT 143.54 281.48 144.64 281.64 ;
      RECT 143.54 281.08 143.7 281.64 ;
      RECT 143.54 281.08 144.64 281.24 ;
      RECT 143.54 282.88 144.64 283.04 ;
      RECT 143.54 282.48 143.7 283.04 ;
      RECT 143.54 282.48 144.64 282.64 ;
      RECT 143.54 284.88 144.64 285.04 ;
      RECT 143.54 284.48 143.7 285.04 ;
      RECT 143.54 284.48 144.64 284.64 ;
      RECT 143.54 286.28 144.64 286.44 ;
      RECT 143.54 285.88 143.7 286.44 ;
      RECT 143.54 285.88 144.64 286.04 ;
      RECT 143.54 288.28 144.64 288.44 ;
      RECT 143.54 287.88 143.7 288.44 ;
      RECT 143.54 287.88 144.64 288.04 ;
      RECT 143.54 289.68 144.64 289.84 ;
      RECT 143.54 289.28 143.7 289.84 ;
      RECT 143.54 289.28 144.64 289.44 ;
      RECT 143.54 291.68 144.64 291.84 ;
      RECT 143.54 291.28 143.7 291.84 ;
      RECT 143.54 291.28 144.64 291.44 ;
      RECT 143.54 293.08 144.64 293.24 ;
      RECT 143.54 292.68 143.7 293.24 ;
      RECT 143.54 292.68 144.64 292.84 ;
      RECT 143.54 295.08 144.64 295.24 ;
      RECT 143.54 294.68 143.7 295.24 ;
      RECT 143.54 294.68 144.64 294.84 ;
      RECT 143.54 296.48 144.64 296.64 ;
      RECT 143.54 296.08 143.7 296.64 ;
      RECT 143.54 296.08 144.64 296.24 ;
      RECT 143.54 298.48 144.64 298.64 ;
      RECT 143.54 298.08 143.7 298.64 ;
      RECT 143.54 298.08 144.64 298.24 ;
      RECT 143.54 299.88 144.64 300.04 ;
      RECT 143.54 299.48 143.7 300.04 ;
      RECT 143.54 299.48 144.64 299.64 ;
      RECT 143.54 301.88 144.64 302.04 ;
      RECT 143.54 301.48 143.7 302.04 ;
      RECT 143.54 301.48 144.64 301.64 ;
      RECT 143.54 303.28 144.64 303.44 ;
      RECT 143.54 302.88 143.7 303.44 ;
      RECT 143.54 302.88 144.64 303.04 ;
      RECT 143.54 305.28 144.64 305.44 ;
      RECT 143.54 304.88 143.7 305.44 ;
      RECT 143.54 304.88 144.64 305.04 ;
      RECT 143.54 306.68 144.64 306.84 ;
      RECT 143.54 306.28 143.7 306.84 ;
      RECT 143.54 306.28 144.64 306.44 ;
      RECT 143.54 308.68 144.64 308.84 ;
      RECT 143.54 308.28 143.7 308.84 ;
      RECT 143.54 308.28 144.64 308.44 ;
      RECT 143.54 310.08 144.64 310.24 ;
      RECT 143.54 309.68 143.7 310.24 ;
      RECT 143.54 309.68 144.64 309.84 ;
      RECT 143.54 312.08 144.64 312.24 ;
      RECT 143.54 311.68 143.7 312.24 ;
      RECT 143.54 311.68 144.64 311.84 ;
      RECT 143.54 313.48 144.64 313.64 ;
      RECT 143.54 313.08 143.7 313.64 ;
      RECT 143.54 313.08 144.64 313.24 ;
      RECT 143.54 315.48 144.64 315.64 ;
      RECT 143.54 315.08 143.7 315.64 ;
      RECT 143.54 315.08 144.64 315.24 ;
      RECT 143.54 316.88 144.64 317.04 ;
      RECT 143.54 316.48 143.7 317.04 ;
      RECT 143.54 316.48 144.64 316.64 ;
      RECT 143.54 318.88 144.64 319.04 ;
      RECT 143.54 318.48 143.7 319.04 ;
      RECT 143.54 318.48 144.64 318.64 ;
      RECT 143.54 320.28 144.64 320.44 ;
      RECT 143.54 319.88 143.7 320.44 ;
      RECT 143.54 319.88 144.64 320.04 ;
      RECT 143.54 322.28 144.64 322.44 ;
      RECT 143.54 321.88 143.7 322.44 ;
      RECT 143.54 321.88 144.64 322.04 ;
      RECT 143.54 323.68 144.64 323.84 ;
      RECT 143.54 323.28 143.7 323.84 ;
      RECT 143.54 323.28 144.64 323.44 ;
      RECT 143.54 325.68 144.64 325.84 ;
      RECT 143.54 325.28 143.7 325.84 ;
      RECT 143.54 325.28 144.64 325.44 ;
      RECT 143.54 327.08 144.64 327.24 ;
      RECT 143.54 326.68 143.7 327.24 ;
      RECT 143.54 326.68 144.64 326.84 ;
      RECT 143.54 329.08 144.64 329.24 ;
      RECT 143.54 328.68 143.7 329.24 ;
      RECT 143.54 328.68 144.64 328.84 ;
      RECT 143.54 330.48 144.64 330.64 ;
      RECT 143.54 330.08 143.7 330.64 ;
      RECT 143.54 330.08 144.64 330.24 ;
      RECT 143.54 332.48 144.64 332.64 ;
      RECT 143.54 332.08 143.7 332.64 ;
      RECT 143.54 332.08 144.64 332.24 ;
      RECT 143.54 333.88 144.64 334.04 ;
      RECT 143.54 333.48 143.7 334.04 ;
      RECT 143.54 333.48 144.64 333.64 ;
      RECT 143.54 335.88 144.64 336.04 ;
      RECT 143.54 335.48 143.7 336.04 ;
      RECT 143.54 335.48 144.64 335.64 ;
      RECT 143.54 337.28 144.64 337.44 ;
      RECT 143.54 336.88 143.7 337.44 ;
      RECT 143.54 336.88 144.64 337.04 ;
      RECT 143.54 339.28 144.64 339.44 ;
      RECT 143.54 338.88 143.7 339.44 ;
      RECT 143.54 338.88 144.64 339.04 ;
      RECT 143.54 340.68 144.64 340.84 ;
      RECT 143.54 340.28 143.7 340.84 ;
      RECT 143.54 340.28 144.64 340.44 ;
      RECT 143.54 342.68 144.64 342.84 ;
      RECT 143.54 342.28 143.7 342.84 ;
      RECT 143.54 342.28 144.64 342.44 ;
      RECT 143.54 344.08 144.64 344.24 ;
      RECT 143.54 343.68 143.7 344.24 ;
      RECT 143.54 343.68 144.64 343.84 ;
      RECT 143.54 346.08 144.64 346.24 ;
      RECT 143.54 345.68 143.7 346.24 ;
      RECT 143.54 345.68 144.64 345.84 ;
      RECT 143.54 347.48 144.64 347.64 ;
      RECT 143.54 347.08 143.7 347.64 ;
      RECT 143.54 347.08 144.64 347.24 ;
      RECT 143.54 349.48 144.64 349.64 ;
      RECT 143.54 349.08 143.7 349.64 ;
      RECT 143.54 349.08 144.64 349.24 ;
      RECT 143.54 350.88 144.64 351.04 ;
      RECT 143.54 350.48 143.7 351.04 ;
      RECT 143.54 350.48 144.64 350.64 ;
      RECT 143.54 352.88 144.64 353.04 ;
      RECT 143.54 352.48 143.7 353.04 ;
      RECT 143.54 352.48 144.64 352.64 ;
      RECT 143.54 354.28 144.64 354.44 ;
      RECT 143.54 353.88 143.7 354.44 ;
      RECT 143.54 353.88 144.64 354.04 ;
      RECT 143.54 356.28 144.64 356.44 ;
      RECT 143.54 355.88 143.7 356.44 ;
      RECT 143.54 355.88 144.64 356.04 ;
      RECT 143.54 357.68 144.64 357.84 ;
      RECT 143.54 357.28 143.7 357.84 ;
      RECT 143.54 357.28 144.64 357.44 ;
      RECT 143.54 359.68 144.64 359.84 ;
      RECT 143.54 359.28 143.7 359.84 ;
      RECT 143.54 359.28 144.64 359.44 ;
      RECT 143.54 361.08 144.64 361.24 ;
      RECT 143.54 360.68 143.7 361.24 ;
      RECT 143.54 360.68 144.64 360.84 ;
      RECT 143.54 363.08 144.64 363.24 ;
      RECT 143.54 362.68 143.7 363.24 ;
      RECT 143.54 362.68 144.64 362.84 ;
      RECT 143.54 364.48 144.64 364.64 ;
      RECT 143.54 364.08 143.7 364.64 ;
      RECT 143.54 364.08 144.64 364.24 ;
      RECT 143.54 366.48 144.64 366.64 ;
      RECT 143.54 366.08 143.7 366.64 ;
      RECT 143.54 366.08 144.64 366.24 ;
      RECT 143.54 367.88 144.64 368.04 ;
      RECT 143.54 367.48 143.7 368.04 ;
      RECT 143.54 367.48 144.64 367.64 ;
      RECT 143.54 369.88 144.64 370.04 ;
      RECT 143.54 369.48 143.7 370.04 ;
      RECT 143.54 369.48 144.64 369.64 ;
      RECT 143.54 371.28 144.64 371.44 ;
      RECT 143.54 370.88 143.7 371.44 ;
      RECT 143.54 370.88 144.64 371.04 ;
      RECT 143.54 373.28 144.64 373.44 ;
      RECT 143.54 372.88 143.7 373.44 ;
      RECT 143.54 372.88 144.64 373.04 ;
      RECT 143.54 374.68 144.64 374.84 ;
      RECT 143.54 374.28 143.7 374.84 ;
      RECT 143.54 374.28 144.64 374.44 ;
      RECT 143.54 376.68 144.64 376.84 ;
      RECT 143.54 376.28 143.7 376.84 ;
      RECT 143.54 376.28 144.64 376.44 ;
      RECT 143.54 378.08 144.64 378.24 ;
      RECT 143.54 377.68 143.7 378.24 ;
      RECT 143.54 377.68 144.64 377.84 ;
      RECT 143.54 380.08 144.64 380.24 ;
      RECT 143.54 379.68 143.7 380.24 ;
      RECT 143.54 379.68 144.64 379.84 ;
      RECT 143.54 381.48 144.64 381.64 ;
      RECT 143.54 381.08 143.7 381.64 ;
      RECT 143.54 381.08 144.64 381.24 ;
      RECT 143.54 383.48 144.64 383.64 ;
      RECT 143.54 383.08 143.7 383.64 ;
      RECT 143.54 383.08 144.64 383.24 ;
      RECT 143.54 384.88 144.64 385.04 ;
      RECT 143.54 384.48 143.7 385.04 ;
      RECT 143.54 384.48 144.64 384.64 ;
      RECT 143.54 386.88 144.64 387.04 ;
      RECT 143.54 386.48 143.7 387.04 ;
      RECT 143.54 386.48 144.64 386.64 ;
      RECT 143.54 388.28 144.64 388.44 ;
      RECT 143.54 387.88 143.7 388.44 ;
      RECT 143.54 387.88 144.64 388.04 ;
      RECT 143.54 390.28 144.64 390.44 ;
      RECT 143.54 389.88 143.7 390.44 ;
      RECT 143.54 389.88 144.64 390.04 ;
      RECT 143.54 391.68 144.64 391.84 ;
      RECT 143.54 391.28 143.7 391.84 ;
      RECT 143.54 391.28 144.64 391.44 ;
      RECT 143.54 393.68 144.64 393.84 ;
      RECT 143.54 393.28 143.7 393.84 ;
      RECT 143.54 393.28 144.64 393.44 ;
      RECT 143.54 395.08 144.64 395.24 ;
      RECT 143.54 394.68 143.7 395.24 ;
      RECT 143.54 394.68 144.64 394.84 ;
      RECT 143.54 397.08 144.64 397.24 ;
      RECT 143.54 396.68 143.7 397.24 ;
      RECT 143.54 396.68 144.64 396.84 ;
      RECT 143.54 398.48 144.64 398.64 ;
      RECT 143.54 398.08 143.7 398.64 ;
      RECT 143.54 398.08 144.64 398.24 ;
      RECT 143.54 400.48 144.64 400.64 ;
      RECT 143.54 400.08 143.7 400.64 ;
      RECT 143.54 400.08 144.64 400.24 ;
      RECT 143.54 401.88 144.64 402.04 ;
      RECT 143.54 401.48 143.7 402.04 ;
      RECT 143.54 401.48 144.64 401.64 ;
      RECT 143.54 403.88 144.64 404.04 ;
      RECT 143.54 403.48 143.7 404.04 ;
      RECT 143.54 403.48 144.64 403.64 ;
      RECT 143.54 405.28 144.64 405.44 ;
      RECT 143.54 404.88 143.7 405.44 ;
      RECT 143.54 404.88 144.64 405.04 ;
      RECT 143.54 407.28 144.64 407.44 ;
      RECT 143.54 406.88 143.7 407.44 ;
      RECT 143.54 406.88 144.64 407.04 ;
      RECT 143.54 408.68 144.64 408.84 ;
      RECT 143.54 408.28 143.7 408.84 ;
      RECT 143.54 408.28 144.64 408.44 ;
      RECT 143.54 410.68 144.64 410.84 ;
      RECT 143.54 410.28 143.7 410.84 ;
      RECT 143.54 410.28 144.64 410.44 ;
      RECT 143.54 412.08 144.64 412.24 ;
      RECT 143.54 411.68 143.7 412.24 ;
      RECT 143.54 411.68 144.64 411.84 ;
      RECT 143.54 414.08 144.64 414.24 ;
      RECT 143.54 413.68 143.7 414.24 ;
      RECT 143.54 413.68 144.64 413.84 ;
      RECT 143.54 415.48 144.64 415.64 ;
      RECT 143.54 415.08 143.7 415.64 ;
      RECT 143.54 415.08 144.64 415.24 ;
      RECT 143.54 417.48 144.64 417.64 ;
      RECT 143.54 417.08 143.7 417.64 ;
      RECT 143.54 417.08 144.64 417.24 ;
      RECT 143.54 418.88 144.64 419.04 ;
      RECT 143.54 418.48 143.7 419.04 ;
      RECT 143.54 418.48 144.64 418.64 ;
      RECT 143.54 420.88 144.64 421.04 ;
      RECT 143.54 420.48 143.7 421.04 ;
      RECT 143.54 420.48 144.64 420.64 ;
      RECT 143.54 422.28 144.64 422.44 ;
      RECT 143.54 421.88 143.7 422.44 ;
      RECT 143.54 421.88 144.64 422.04 ;
      RECT 143.54 424.28 144.64 424.44 ;
      RECT 143.54 423.88 143.7 424.44 ;
      RECT 143.54 423.88 144.64 424.04 ;
      RECT 143.54 425.68 144.64 425.84 ;
      RECT 143.54 425.28 143.7 425.84 ;
      RECT 143.54 425.28 144.64 425.44 ;
      RECT 143.54 427.68 144.64 427.84 ;
      RECT 143.54 427.28 143.7 427.84 ;
      RECT 143.54 427.28 144.64 427.44 ;
      RECT 143.54 429.08 144.64 429.24 ;
      RECT 143.54 428.68 143.7 429.24 ;
      RECT 143.54 428.68 144.64 428.84 ;
      RECT 143.54 431.08 144.64 431.24 ;
      RECT 143.54 430.68 143.7 431.24 ;
      RECT 143.54 430.68 144.64 430.84 ;
      RECT 143.54 432.48 144.64 432.64 ;
      RECT 143.54 432.08 143.7 432.64 ;
      RECT 143.54 432.08 144.64 432.24 ;
      RECT 143.54 434.48 144.64 434.64 ;
      RECT 143.54 434.08 143.7 434.64 ;
      RECT 143.54 434.08 144.64 434.24 ;
      RECT 143.54 435.88 144.64 436.04 ;
      RECT 143.54 435.48 143.7 436.04 ;
      RECT 143.54 435.48 144.64 435.64 ;
      RECT 143.54 437.88 144.64 438.04 ;
      RECT 143.54 437.48 143.7 438.04 ;
      RECT 143.54 437.48 144.64 437.64 ;
      RECT 143.54 439.28 144.64 439.44 ;
      RECT 143.54 438.88 143.7 439.44 ;
      RECT 143.54 438.88 144.64 439.04 ;
      RECT 143.54 441.28 144.64 441.44 ;
      RECT 143.54 440.88 143.7 441.44 ;
      RECT 143.54 440.88 144.64 441.04 ;
      RECT 143.54 442.68 144.64 442.84 ;
      RECT 143.54 442.28 143.7 442.84 ;
      RECT 143.54 442.28 144.64 442.44 ;
      RECT 143.54 444.68 144.64 444.84 ;
      RECT 143.54 444.28 143.7 444.84 ;
      RECT 143.54 444.28 144.64 444.44 ;
      RECT 143.54 446.08 144.64 446.24 ;
      RECT 143.54 445.68 143.7 446.24 ;
      RECT 143.54 445.68 144.64 445.84 ;
      RECT 143.54 448.08 144.64 448.24 ;
      RECT 143.54 447.68 143.7 448.24 ;
      RECT 143.54 447.68 144.64 447.84 ;
      RECT 143.54 449.48 144.64 449.64 ;
      RECT 143.54 449.08 143.7 449.64 ;
      RECT 143.54 449.08 144.64 449.24 ;
      RECT 143.54 451.48 144.64 451.64 ;
      RECT 143.54 451.08 143.7 451.64 ;
      RECT 143.54 451.08 144.64 451.24 ;
      RECT 143.54 452.88 144.64 453.04 ;
      RECT 143.54 452.48 143.7 453.04 ;
      RECT 143.54 452.48 144.64 452.64 ;
      RECT 143.54 454.88 144.64 455.04 ;
      RECT 143.54 454.48 143.7 455.04 ;
      RECT 143.54 454.48 144.64 454.64 ;
      RECT 143.54 456.28 144.64 456.44 ;
      RECT 143.54 455.88 143.7 456.44 ;
      RECT 143.54 455.88 144.64 456.04 ;
      RECT 143.54 458.28 144.64 458.44 ;
      RECT 143.54 457.88 143.7 458.44 ;
      RECT 143.54 457.88 144.64 458.04 ;
      RECT 143.54 459.68 144.64 459.84 ;
      RECT 143.54 459.28 143.7 459.84 ;
      RECT 143.54 459.28 144.64 459.44 ;
      RECT 143.54 461.68 144.64 461.84 ;
      RECT 143.54 461.28 143.7 461.84 ;
      RECT 143.54 461.28 144.64 461.44 ;
      RECT 143.54 463.08 144.64 463.24 ;
      RECT 143.54 462.68 143.7 463.24 ;
      RECT 143.54 462.68 144.64 462.84 ;
      RECT 143.54 465.08 144.64 465.24 ;
      RECT 143.54 464.68 143.7 465.24 ;
      RECT 143.54 464.68 144.64 464.84 ;
      RECT 143.54 466.48 144.64 466.64 ;
      RECT 143.54 466.08 143.7 466.64 ;
      RECT 143.54 466.08 144.64 466.24 ;
      RECT 143.54 468.48 144.64 468.64 ;
      RECT 143.54 468.08 143.7 468.64 ;
      RECT 143.54 468.08 144.64 468.24 ;
      RECT 143.54 469.88 144.64 470.04 ;
      RECT 143.54 469.48 143.7 470.04 ;
      RECT 143.54 469.48 144.64 469.64 ;
      RECT 143.54 471.88 144.64 472.04 ;
      RECT 143.54 471.48 143.7 472.04 ;
      RECT 143.54 471.48 144.64 471.64 ;
      RECT 143.54 473.28 144.64 473.44 ;
      RECT 143.54 472.88 143.7 473.44 ;
      RECT 143.54 472.88 144.64 473.04 ;
      RECT 143.54 475.28 144.64 475.44 ;
      RECT 143.54 474.88 143.7 475.44 ;
      RECT 143.54 474.88 144.64 475.04 ;
      RECT 143.54 476.68 144.64 476.84 ;
      RECT 143.54 476.28 143.7 476.84 ;
      RECT 143.54 476.28 144.64 476.44 ;
      RECT 143.54 478.68 144.64 478.84 ;
      RECT 143.54 478.28 143.7 478.84 ;
      RECT 143.54 478.28 144.64 478.44 ;
      RECT 143.54 480.08 144.64 480.24 ;
      RECT 143.54 479.68 143.7 480.24 ;
      RECT 143.54 479.68 144.64 479.84 ;
      RECT 143.54 482.08 144.64 482.24 ;
      RECT 143.54 481.68 143.7 482.24 ;
      RECT 143.54 481.68 144.64 481.84 ;
      RECT 143.54 483.48 144.64 483.64 ;
      RECT 143.54 483.08 143.7 483.64 ;
      RECT 143.54 483.08 144.64 483.24 ;
      RECT 143.54 485.48 144.64 485.64 ;
      RECT 143.54 485.08 143.7 485.64 ;
      RECT 143.54 485.08 144.64 485.24 ;
      RECT 143.54 486.88 144.64 487.04 ;
      RECT 143.54 486.48 143.7 487.04 ;
      RECT 143.54 486.48 144.64 486.64 ;
      RECT 143.54 488.88 144.64 489.04 ;
      RECT 143.54 488.48 143.7 489.04 ;
      RECT 143.54 488.48 144.64 488.64 ;
      RECT 143.54 490.28 144.64 490.44 ;
      RECT 143.54 489.88 143.7 490.44 ;
      RECT 143.54 489.88 144.64 490.04 ;
      RECT 143.54 492.28 144.64 492.44 ;
      RECT 143.54 491.88 143.7 492.44 ;
      RECT 143.54 491.88 144.64 492.04 ;
      RECT 143.54 493.68 144.64 493.84 ;
      RECT 143.54 493.28 143.7 493.84 ;
      RECT 143.54 493.28 144.64 493.44 ;
      RECT 143.54 495.68 144.64 495.84 ;
      RECT 143.54 495.28 143.7 495.84 ;
      RECT 143.54 495.28 144.64 495.44 ;
      RECT 143.54 497.08 144.64 497.24 ;
      RECT 143.54 496.68 143.7 497.24 ;
      RECT 143.54 496.68 144.64 496.84 ;
      RECT 143.54 499.08 144.64 499.24 ;
      RECT 143.54 498.68 143.7 499.24 ;
      RECT 143.54 498.68 144.64 498.84 ;
      RECT 143.54 500.48 144.64 500.64 ;
      RECT 143.54 500.08 143.7 500.64 ;
      RECT 143.54 500.08 144.64 500.24 ;
      RECT 143.54 502.48 144.64 502.64 ;
      RECT 143.54 502.08 143.7 502.64 ;
      RECT 143.54 502.08 144.64 502.24 ;
      RECT 143.54 503.88 144.64 504.04 ;
      RECT 143.54 503.48 143.7 504.04 ;
      RECT 143.54 503.48 144.64 503.64 ;
      RECT 144.38 30.98 144.54 32.25 ;
      RECT 144.35 29.19 144.51 31.14 ;
      RECT 143.6 29.87 144.51 30.11 ;
      RECT 144.27 28.58 144.43 29.37 ;
      RECT 143.35 37.35 144.43 37.51 ;
      RECT 144.27 35.68 144.43 37.51 ;
      RECT 143.31 35.68 143.47 36.68 ;
      RECT 143.21 35.68 144.53 35.84 ;
      RECT 144.37 34.58 144.53 35.84 ;
      RECT 143.21 34.58 143.37 35.84 ;
      RECT 144.27 34.58 144.53 34.86 ;
      RECT 143.21 34.58 143.47 34.86 ;
      RECT 143.79 42.53 143.95 46.23 ;
      RECT 143.31 42.53 144.43 42.69 ;
      RECT 144.27 37.99 144.43 42.69 ;
      RECT 143.31 37.99 143.47 42.69 ;
      RECT 143.31 43.34 143.47 47.95 ;
      RECT 143.31 46.47 144.43 46.63 ;
      RECT 144.27 43.34 144.43 46.63 ;
      RECT 143.53 51.95 144.21 52.11 ;
      RECT 143.79 51.6 143.95 52.11 ;
      RECT 142.94 29.34 143.1 32.11 ;
      RECT 142.94 29.55 144.19 29.71 ;
      RECT 142.94 29.34 143.23 29.71 ;
      RECT 141.86 29.34 143.23 29.5 ;
      RECT 142.82 29.06 142.98 29.5 ;
      RECT 141.86 29.06 142.02 29.5 ;
      RECT 142.13 22.69 142.29 23.27 ;
      RECT 142.13 22.69 142.93 22.85 ;
      RECT 142.77 21.55 142.93 22.85 ;
      RECT 142.77 21.55 144.03 21.71 ;
      RECT 135.81 505.64 143.38 505.8 ;
      RECT 131.44 505.64 135.26 505.8 ;
      RECT 135.1 504.68 135.26 505.8 ;
      RECT 135.81 504.68 135.97 505.8 ;
      RECT 130.68 504.68 143.97 504.84 ;
      RECT 143.79 28.09 143.95 29.37 ;
      RECT 143.27 28.09 143.95 28.32 ;
      RECT 143.79 47.16 143.95 51.33 ;
      RECT 141.87 47.16 142.03 51.33 ;
      RECT 141.87 48.4 143.95 48.59 ;
      RECT 142.83 47.14 142.99 48.59 ;
      RECT 143.33 42.85 143.63 43.09 ;
      RECT 143.05 42.85 143.63 43.03 ;
      RECT 143.08 6.24 143.36 7.12 ;
      RECT 142.62 6.24 143.57 6.84 ;
      RECT 142.34 28.22 142.5 29.18 ;
      RECT 142.34 28.22 143.01 28.38 ;
      RECT 142.85 28.1 143.01 28.38 ;
      RECT 142.75 509.04 142.91 509.54 ;
      RECT 141.77 509.04 141.93 509.54 ;
      RECT 141.77 509.04 142.91 509.2 ;
      RECT 142.26 507.6 142.42 509.2 ;
      RECT 141.77 507.6 142.91 507.76 ;
      RECT 142.75 507.26 142.91 507.76 ;
      RECT 141.77 507.26 141.93 507.76 ;
      RECT 141.96 30.5 142.78 30.66 ;
      RECT 142.62 30.29 142.78 30.66 ;
      RECT 142.19 42.85 142.49 43.09 ;
      RECT 142.19 42.85 142.77 43.03 ;
      RECT 141.23 52.33 142.67 52.55 ;
      RECT 142.45 51.48 142.67 52.55 ;
      RECT 141.23 51.44 141.45 52.55 ;
      RECT 142.35 48.78 142.51 51.77 ;
      RECT 141.39 46.79 141.55 51.77 ;
      RECT 141.39 46.79 142.19 47 ;
      RECT 140.91 46.79 142.19 46.96 ;
      RECT 140.91 43.19 141.07 46.96 ;
      RECT 141.39 37.35 142.47 37.51 ;
      RECT 141.39 35.68 141.55 37.51 ;
      RECT 142.35 35.68 142.51 36.68 ;
      RECT 141.29 35.68 142.61 35.84 ;
      RECT 142.45 34.58 142.61 35.84 ;
      RECT 141.29 34.58 141.45 35.84 ;
      RECT 142.35 34.58 142.61 34.86 ;
      RECT 141.29 34.58 141.55 34.86 ;
      RECT 141.87 42.53 142.03 46.23 ;
      RECT 141.39 42.53 142.51 42.69 ;
      RECT 142.35 37.99 142.51 42.69 ;
      RECT 141.39 37.99 141.55 42.69 ;
      RECT 142.35 43.34 142.51 47.95 ;
      RECT 141.39 46.47 142.51 46.63 ;
      RECT 141.39 43.34 141.55 46.63 ;
      RECT 141.82 32.74 142.34 32.9 ;
      RECT 141.82 30.84 141.98 32.9 ;
      RECT 141.61 51.95 142.29 52.11 ;
      RECT 141.87 51.6 142.03 52.11 ;
      RECT 141.41 42.85 141.71 43.09 ;
      RECT 141.13 42.85 141.71 43.03 ;
      RECT 141.01 509.04 141.17 509.54 ;
      RECT 140.03 509.04 140.19 509.54 ;
      RECT 140.03 509.04 141.17 509.2 ;
      RECT 140.52 507.6 140.68 509.2 ;
      RECT 140.03 507.6 141.17 507.76 ;
      RECT 141.01 507.26 141.17 507.76 ;
      RECT 140.03 507.26 140.19 507.76 ;
      RECT 138.39 12.34 138.67 12.62 ;
      RECT 137.47 12.34 137.75 12.62 ;
      RECT 135.07 12.34 135.35 12.62 ;
      RECT 134.15 12.34 134.43 12.62 ;
      RECT 131.59 12.34 131.87 12.62 ;
      RECT 130.67 12.34 130.95 12.62 ;
      RECT 128.27 12.34 128.55 12.62 ;
      RECT 127.35 12.34 127.63 12.62 ;
      RECT 138.51 11.75 138.67 12.62 ;
      RECT 137.47 11.75 137.63 12.62 ;
      RECT 135.19 11.75 135.35 12.62 ;
      RECT 134.15 11.75 134.31 12.62 ;
      RECT 131.71 11.75 131.87 12.62 ;
      RECT 130.67 11.75 130.83 12.62 ;
      RECT 128.39 11.75 128.55 12.62 ;
      RECT 127.35 11.75 127.51 12.62 ;
      RECT 139.73 8.38 139.89 12.03 ;
      RECT 138.63 9.02 138.79 12.03 ;
      RECT 137.43 9.02 137.59 12.03 ;
      RECT 136.33 8.38 136.49 12.03 ;
      RECT 135.23 9.02 135.39 12.03 ;
      RECT 134.03 9.02 134.19 12.03 ;
      RECT 132.93 8.38 133.09 12.03 ;
      RECT 131.83 9.02 131.99 12.03 ;
      RECT 130.63 9.02 130.79 12.03 ;
      RECT 129.53 8.38 129.69 12.03 ;
      RECT 128.43 9.02 128.59 12.03 ;
      RECT 127.23 9.02 127.39 12.03 ;
      RECT 126.13 8.38 126.29 12.03 ;
      RECT 126.13 9.02 139.89 9.3 ;
      RECT 139.05 8.38 139.29 9.3 ;
      RECT 138.36 8.38 138.6 9.3 ;
      RECT 137.61 8.38 137.85 9.3 ;
      RECT 136.93 8.38 137.17 9.3 ;
      RECT 135.65 8.38 135.89 9.3 ;
      RECT 134.97 8.38 135.21 9.3 ;
      RECT 134.22 8.38 134.46 9.3 ;
      RECT 133.53 8.38 133.77 9.3 ;
      RECT 132.25 8.38 132.49 9.3 ;
      RECT 131.56 8.38 131.8 9.3 ;
      RECT 130.81 8.38 131.05 9.3 ;
      RECT 130.13 8.38 130.37 9.3 ;
      RECT 128.85 8.38 129.09 9.3 ;
      RECT 128.17 8.38 128.41 9.3 ;
      RECT 127.42 8.38 127.66 9.3 ;
      RECT 126.73 8.38 126.97 9.3 ;
      RECT 139.73 17.6 139.89 23.81 ;
      RECT 139.25 22.38 139.89 22.54 ;
      RECT 139.31 27.37 139.47 31.49 ;
      RECT 139.31 27.37 139.89 27.53 ;
      RECT 139.73 24.64 139.89 27.53 ;
      RECT 139.73 54.16 139.89 57.42 ;
      RECT 139.31 54.16 139.89 54.88 ;
      RECT 139.31 50.8 139.47 54.88 ;
      RECT 139.73 58.24 139.89 64 ;
      RECT 139.25 59.51 139.89 59.67 ;
      RECT 88.73 67.14 139.89 67.3 ;
      RECT 139.41 64.6 139.89 67.3 ;
      RECT 138.51 65.19 138.67 67.3 ;
      RECT 137.55 65.19 137.71 67.3 ;
      RECT 136.01 64.6 136.81 67.3 ;
      RECT 136.65 63.97 136.81 67.3 ;
      RECT 135.11 65.19 135.27 67.3 ;
      RECT 134.15 65.19 134.31 67.3 ;
      RECT 132.61 64.6 133.41 67.3 ;
      RECT 133.25 63.96 133.41 67.3 ;
      RECT 131.71 65.19 131.87 67.3 ;
      RECT 130.75 65.19 130.91 67.3 ;
      RECT 129.21 64.6 130.01 67.3 ;
      RECT 129.85 63.97 130.01 67.3 ;
      RECT 128.31 65.19 128.47 67.3 ;
      RECT 127.35 65.19 127.51 67.3 ;
      RECT 125.81 64.6 126.61 67.3 ;
      RECT 126.45 63.96 126.61 67.3 ;
      RECT 124.91 65.19 125.07 67.3 ;
      RECT 123.95 65.19 124.11 67.3 ;
      RECT 122.41 64.6 123.21 67.3 ;
      RECT 123.05 63.97 123.21 67.3 ;
      RECT 121.51 65.19 121.67 67.3 ;
      RECT 120.55 65.19 120.71 67.3 ;
      RECT 119.01 64.6 119.81 67.3 ;
      RECT 119.65 63.96 119.81 67.3 ;
      RECT 118.11 65.19 118.27 67.3 ;
      RECT 117.15 65.19 117.31 67.3 ;
      RECT 115.61 64.6 116.41 67.3 ;
      RECT 116.25 63.97 116.41 67.3 ;
      RECT 114.71 65.19 114.87 67.3 ;
      RECT 113.75 65.19 113.91 67.3 ;
      RECT 112.21 64.6 113.01 67.3 ;
      RECT 112.85 63.96 113.01 67.3 ;
      RECT 111.31 65.19 111.47 67.3 ;
      RECT 110.35 65.19 110.51 67.3 ;
      RECT 108.81 64.6 109.61 67.3 ;
      RECT 109.45 63.97 109.61 67.3 ;
      RECT 107.91 65.19 108.07 67.3 ;
      RECT 106.95 65.19 107.11 67.3 ;
      RECT 105.41 64.6 106.21 67.3 ;
      RECT 106.05 63.96 106.21 67.3 ;
      RECT 104.51 65.19 104.67 67.3 ;
      RECT 103.55 65.19 103.71 67.3 ;
      RECT 102.01 64.6 102.81 67.3 ;
      RECT 102.65 63.97 102.81 67.3 ;
      RECT 101.11 65.19 101.27 67.3 ;
      RECT 100.15 65.19 100.31 67.3 ;
      RECT 98.61 64.6 99.41 67.3 ;
      RECT 99.25 63.96 99.41 67.3 ;
      RECT 97.71 65.19 97.87 67.3 ;
      RECT 96.75 65.19 96.91 67.3 ;
      RECT 95.21 64.6 96.01 67.3 ;
      RECT 95.85 63.97 96.01 67.3 ;
      RECT 94.31 65.19 94.47 67.3 ;
      RECT 93.35 65.19 93.51 67.3 ;
      RECT 91.81 64.6 92.61 67.3 ;
      RECT 92.45 63.96 92.61 67.3 ;
      RECT 90.91 65.19 91.07 67.3 ;
      RECT 89.95 65.19 90.11 67.3 ;
      RECT 88.73 64.6 89.21 67.3 ;
      RECT 89.05 63.97 89.21 67.3 ;
      RECT 139.41 63.96 139.57 67.3 ;
      RECT 136.01 63.97 136.17 67.3 ;
      RECT 132.61 63.96 132.77 67.3 ;
      RECT 129.21 63.97 129.37 67.3 ;
      RECT 125.81 63.96 125.97 67.3 ;
      RECT 122.41 63.97 122.57 67.3 ;
      RECT 119.01 63.96 119.17 67.3 ;
      RECT 115.61 63.97 115.77 67.3 ;
      RECT 112.21 63.96 112.37 67.3 ;
      RECT 108.81 63.97 108.97 67.3 ;
      RECT 105.41 63.96 105.57 67.3 ;
      RECT 102.01 63.97 102.17 67.3 ;
      RECT 98.61 63.96 98.77 67.3 ;
      RECT 95.21 63.97 95.37 67.3 ;
      RECT 91.81 63.96 91.97 67.3 ;
      RECT 137.57 55.09 138.83 55.25 ;
      RECT 138.67 49.77 138.83 55.25 ;
      RECT 138.67 49.77 139.55 49.93 ;
      RECT 139.39 32.48 139.55 49.93 ;
      RECT 138.73 45.9 139.55 46.06 ;
      RECT 138.73 36.23 139.55 36.39 ;
      RECT 138.67 32.48 139.55 32.64 ;
      RECT 138.67 27.04 138.83 32.64 ;
      RECT 137.57 27.04 138.83 27.2 ;
      RECT 137.47 26.46 139.49 26.62 ;
      RECT 139.33 25.35 139.49 26.62 ;
      RECT 139.25 22.91 139.41 25.51 ;
      RECT 139.25 56.46 139.41 59.14 ;
      RECT 139.33 55.49 139.49 56.62 ;
      RECT 137.47 55.49 139.49 55.65 ;
      RECT 139.27 509.04 139.43 509.54 ;
      RECT 138.29 509.04 138.45 509.54 ;
      RECT 138.29 509.04 139.43 509.2 ;
      RECT 138.78 507.6 138.94 509.2 ;
      RECT 138.29 507.6 139.43 507.76 ;
      RECT 139.27 507.26 139.43 507.76 ;
      RECT 138.29 507.25 138.45 507.76 ;
      RECT 138.93 25.79 139.17 26.07 ;
      RECT 138.93 21.94 139.09 26.07 ;
      RECT 138.93 21.94 139.21 22.18 ;
      RECT 138.99 15.28 139.15 22.18 ;
      RECT 138.03 15.28 138.19 20.88 ;
      RECT 137.07 15.28 137.23 20.88 ;
      RECT 137.07 17.14 139.15 17.3 ;
      RECT 138.99 59.87 139.15 66.77 ;
      RECT 138.03 61.17 138.19 66.77 ;
      RECT 137.07 61.17 137.23 66.77 ;
      RECT 137.07 64.75 139.15 64.91 ;
      RECT 138.93 59.87 139.21 60.11 ;
      RECT 138.93 56.02 139.09 60.11 ;
      RECT 138.93 56.02 139.17 56.3 ;
      RECT 137.07 35.91 139.15 36.07 ;
      RECT 138.99 32.85 139.15 36.07 ;
      RECT 138.03 27.43 138.19 36.07 ;
      RECT 137.07 32.85 137.23 36.07 ;
      RECT 137.13 27.43 138.19 27.59 ;
      RECT 137.13 23.41 137.29 27.59 ;
      RECT 137.13 26.14 138.29 26.3 ;
      RECT 138.13 25.01 138.29 26.3 ;
      RECT 137.13 25 137.33 26.3 ;
      RECT 138.13 21.38 138.29 23.81 ;
      RECT 137.17 21.38 137.33 23.55 ;
      RECT 137.17 21.38 138.29 21.54 ;
      RECT 137.17 60.51 138.29 60.67 ;
      RECT 138.13 58.24 138.29 60.67 ;
      RECT 137.17 58.5 137.33 60.67 ;
      RECT 137.13 55.81 137.29 58.64 ;
      RECT 138.13 55.81 138.29 57.09 ;
      RECT 137.11 55.81 137.33 57.09 ;
      RECT 137.11 55.81 138.29 55.97 ;
      RECT 137.11 54.64 137.27 57.09 ;
      RECT 137.11 54.64 138.19 54.8 ;
      RECT 138.03 46.22 138.19 54.8 ;
      RECT 138.99 46.22 139.15 49.44 ;
      RECT 137.07 46.22 137.23 49.44 ;
      RECT 137.07 46.22 139.15 46.38 ;
      RECT 138.43 12.8 139.09 13.06 ;
      RECT 138.85 12.19 139.09 13.06 ;
      RECT 138.91 41.08 139.07 45.17 ;
      RECT 138.75 41.08 139.07 41.24 ;
      RECT 138.61 21.06 138.77 26.28 ;
      RECT 137.65 24.37 137.81 25.98 ;
      RECT 137.45 24.37 138.77 24.53 ;
      RECT 137.45 23.67 137.61 24.53 ;
      RECT 137.45 23.67 137.81 23.83 ;
      RECT 137.65 21.7 137.81 23.83 ;
      RECT 136.95 21.06 138.83 21.22 ;
      RECT 136.95 60.83 138.83 60.99 ;
      RECT 138.61 55.81 138.77 60.99 ;
      RECT 137.65 58.22 137.81 60.35 ;
      RECT 137.45 58.22 137.81 58.38 ;
      RECT 137.45 57.25 137.61 58.38 ;
      RECT 137.45 57.25 138.77 57.41 ;
      RECT 137.65 56.13 137.81 57.41 ;
      RECT 138.51 14.52 138.67 16.86 ;
      RECT 138.64 13.22 138.8 14.84 ;
      RECT 138.51 32.85 138.67 35.75 ;
      RECT 138.35 31.09 138.51 33.01 ;
      RECT 138.35 49.44 138.51 51.3 ;
      RECT 138.51 46.54 138.67 49.6 ;
      RECT 138.43 38.57 138.59 45.17 ;
      RECT 138.13 38.57 138.59 38.73 ;
      RECT 138.13 36.23 138.29 38.73 ;
      RECT 137.77 36.23 138.45 36.39 ;
      RECT 137.65 45.9 138.45 46.06 ;
      RECT 137.65 44.89 137.81 46.06 ;
      RECT 137.63 38.57 137.79 45.17 ;
      RECT 138.03 10.09 138.19 14.2 ;
      RECT 137.13 12.9 138.19 13.06 ;
      RECT 137.13 12.19 137.29 13.06 ;
      RECT 137.55 14.52 137.71 16.86 ;
      RECT 137.42 13.22 137.58 14.84 ;
      RECT 137.55 31.09 137.71 35.75 ;
      RECT 137.45 32.25 137.71 32.53 ;
      RECT 137.51 49.75 137.71 51.3 ;
      RECT 137.55 46.54 137.71 51.3 ;
      RECT 137.53 509.04 137.69 509.54 ;
      RECT 137.04 509.04 137.69 509.2 ;
      RECT 137.04 507.6 137.2 509.2 ;
      RECT 137.04 507.6 137.69 507.76 ;
      RECT 137.53 507.25 137.69 507.76 ;
      RECT 137.11 49.6 137.27 51.7 ;
      RECT 136.67 49.6 137.27 49.76 ;
      RECT 136.67 32.06 136.83 49.76 ;
      RECT 136.67 45.9 137.49 46.06 ;
      RECT 136.67 36.23 137.49 36.39 ;
      RECT 136.67 32.06 137.27 32.22 ;
      RECT 137.11 30.54 137.27 32.22 ;
      RECT 137.15 41.08 137.31 45.17 ;
      RECT 137.15 41.08 137.47 41.24 ;
      RECT 136.33 31.49 136.49 32.02 ;
      RECT 135.87 31.49 136.95 31.65 ;
      RECT 136.79 27.38 136.95 31.65 ;
      RECT 135.87 27.38 136.03 31.65 ;
      RECT 135.87 27.38 136.95 27.54 ;
      RECT 136.33 26.91 136.49 27.54 ;
      RECT 135.87 51.06 136.95 55.29 ;
      RECT 136.33 50.27 136.49 55.29 ;
      RECT 136.69 49.92 136.85 50.9 ;
      RECT 135.97 49.92 136.13 50.9 ;
      RECT 135.97 49.92 136.85 50.08 ;
      RECT 136.33 45.65 136.49 50.08 ;
      RECT 135.55 49.6 135.71 51.7 ;
      RECT 135.55 49.6 136.15 49.76 ;
      RECT 135.99 32.06 136.15 49.76 ;
      RECT 135.33 45.9 136.15 46.06 ;
      RECT 135.33 36.23 136.15 36.39 ;
      RECT 135.55 32.06 136.15 32.22 ;
      RECT 135.55 30.54 135.71 32.22 ;
      RECT 134.05 21.06 134.21 26.28 ;
      RECT 135.01 24.37 135.17 25.98 ;
      RECT 134.05 24.37 135.37 24.53 ;
      RECT 135.21 23.67 135.37 24.53 ;
      RECT 135.01 23.67 135.37 23.83 ;
      RECT 135.01 21.7 135.17 23.83 ;
      RECT 133.99 21.06 135.87 21.22 ;
      RECT 133.99 60.83 135.87 60.99 ;
      RECT 134.05 55.81 134.21 60.99 ;
      RECT 135.01 58.22 135.17 60.35 ;
      RECT 135.01 58.22 135.37 58.38 ;
      RECT 135.21 57.25 135.37 58.38 ;
      RECT 134.05 57.25 135.37 57.41 ;
      RECT 135.01 56.13 135.17 57.41 ;
      RECT 133.65 25.79 133.89 26.07 ;
      RECT 133.73 21.94 133.89 26.07 ;
      RECT 133.61 21.94 133.89 22.18 ;
      RECT 133.67 15.28 133.83 22.18 ;
      RECT 135.59 15.28 135.75 20.88 ;
      RECT 134.63 15.28 134.79 20.88 ;
      RECT 133.67 17.14 135.75 17.3 ;
      RECT 133.67 35.91 135.75 36.07 ;
      RECT 135.59 32.85 135.75 36.07 ;
      RECT 134.63 27.43 134.79 36.07 ;
      RECT 133.67 32.85 133.83 36.07 ;
      RECT 134.63 27.43 135.69 27.59 ;
      RECT 135.53 23.41 135.69 27.59 ;
      RECT 134.53 26.14 135.69 26.3 ;
      RECT 135.49 25 135.69 26.3 ;
      RECT 134.53 25.01 134.69 26.3 ;
      RECT 134.53 21.38 134.69 23.81 ;
      RECT 135.49 21.38 135.65 23.55 ;
      RECT 134.53 21.38 135.65 21.54 ;
      RECT 134.53 60.51 135.65 60.67 ;
      RECT 135.49 58.5 135.65 60.67 ;
      RECT 135.53 55.81 135.65 60.67 ;
      RECT 134.53 58.24 134.69 60.67 ;
      RECT 135.55 54.64 135.69 58.64 ;
      RECT 135.49 55.81 135.71 57.09 ;
      RECT 135.55 54.64 135.71 57.09 ;
      RECT 134.53 55.81 134.69 57.09 ;
      RECT 134.53 55.81 135.71 55.97 ;
      RECT 134.63 54.64 135.71 54.8 ;
      RECT 134.63 46.22 134.79 54.8 ;
      RECT 135.59 46.22 135.75 49.44 ;
      RECT 133.67 46.22 133.83 49.44 ;
      RECT 133.67 46.22 135.75 46.38 ;
      RECT 135.59 61.17 135.75 66.77 ;
      RECT 134.63 61.17 134.79 66.77 ;
      RECT 133.67 59.87 133.83 66.77 ;
      RECT 133.67 64.75 135.75 64.91 ;
      RECT 133.61 59.87 133.89 60.11 ;
      RECT 133.73 56.02 133.89 60.11 ;
      RECT 133.65 56.02 133.89 56.3 ;
      RECT 134.63 10.09 134.79 14.2 ;
      RECT 134.63 12.9 135.69 13.06 ;
      RECT 135.53 12.19 135.69 13.06 ;
      RECT 135.51 41.08 135.67 45.17 ;
      RECT 135.35 41.08 135.67 41.24 ;
      RECT 131.12 506.12 134.79 506.28 ;
      RECT 127.66 506.12 129.36 506.28 ;
      RECT 135.49 505.02 135.65 506.12 ;
      RECT 134.63 505.96 135.65 506.12 ;
      RECT 131.12 505.16 131.28 506.28 ;
      RECT 127.66 505.16 127.82 506.28 ;
      RECT 127.66 505.16 134.79 505.32 ;
      RECT 129.08 71 131.27 71.16 ;
      RECT 135.48 69.96 135.64 71.08 ;
      RECT 131.04 70.92 135.64 71.08 ;
      RECT 127.56 70.92 129.36 71.08 ;
      RECT 127.56 69.96 127.72 71.08 ;
      RECT 127.56 69.96 135.64 70.12 ;
      RECT 127.56 72.4 135.64 72.56 ;
      RECT 135.48 71.44 135.64 72.56 ;
      RECT 127.56 71.44 127.72 72.56 ;
      RECT 131.04 71.44 135.64 71.6 ;
      RECT 127.56 71.44 129.36 71.6 ;
      RECT 129.08 71.36 131.27 71.52 ;
      RECT 129.08 74.4 131.27 74.56 ;
      RECT 135.48 73.36 135.64 74.48 ;
      RECT 131.04 74.32 135.64 74.48 ;
      RECT 127.56 74.32 129.36 74.48 ;
      RECT 127.56 73.36 127.72 74.48 ;
      RECT 127.56 73.36 135.64 73.52 ;
      RECT 127.56 75.8 135.64 75.96 ;
      RECT 135.48 74.84 135.64 75.96 ;
      RECT 127.56 74.84 127.72 75.96 ;
      RECT 131.04 74.84 135.64 75 ;
      RECT 127.56 74.84 129.36 75 ;
      RECT 129.08 74.76 131.27 74.92 ;
      RECT 129.08 77.8 131.27 77.96 ;
      RECT 135.48 76.76 135.64 77.88 ;
      RECT 131.04 77.72 135.64 77.88 ;
      RECT 127.56 77.72 129.36 77.88 ;
      RECT 127.56 76.76 127.72 77.88 ;
      RECT 127.56 76.76 135.64 76.92 ;
      RECT 127.56 79.2 135.64 79.36 ;
      RECT 135.48 78.24 135.64 79.36 ;
      RECT 127.56 78.24 127.72 79.36 ;
      RECT 131.04 78.24 135.64 78.4 ;
      RECT 127.56 78.24 129.36 78.4 ;
      RECT 129.08 78.16 131.27 78.32 ;
      RECT 129.08 81.2 131.27 81.36 ;
      RECT 135.48 80.16 135.64 81.28 ;
      RECT 131.04 81.12 135.64 81.28 ;
      RECT 127.56 81.12 129.36 81.28 ;
      RECT 127.56 80.16 127.72 81.28 ;
      RECT 127.56 80.16 135.64 80.32 ;
      RECT 127.56 82.6 135.64 82.76 ;
      RECT 135.48 81.64 135.64 82.76 ;
      RECT 127.56 81.64 127.72 82.76 ;
      RECT 131.04 81.64 135.64 81.8 ;
      RECT 127.56 81.64 129.36 81.8 ;
      RECT 129.08 81.56 131.27 81.72 ;
      RECT 129.08 84.6 131.27 84.76 ;
      RECT 135.48 83.56 135.64 84.68 ;
      RECT 131.04 84.52 135.64 84.68 ;
      RECT 127.56 84.52 129.36 84.68 ;
      RECT 127.56 83.56 127.72 84.68 ;
      RECT 127.56 83.56 135.64 83.72 ;
      RECT 127.56 86 135.64 86.16 ;
      RECT 135.48 85.04 135.64 86.16 ;
      RECT 127.56 85.04 127.72 86.16 ;
      RECT 131.04 85.04 135.64 85.2 ;
      RECT 127.56 85.04 129.36 85.2 ;
      RECT 129.08 84.96 131.27 85.12 ;
      RECT 129.08 88 131.27 88.16 ;
      RECT 135.48 86.96 135.64 88.08 ;
      RECT 131.04 87.92 135.64 88.08 ;
      RECT 127.56 87.92 129.36 88.08 ;
      RECT 127.56 86.96 127.72 88.08 ;
      RECT 127.56 86.96 135.64 87.12 ;
      RECT 127.56 89.4 135.64 89.56 ;
      RECT 135.48 88.44 135.64 89.56 ;
      RECT 127.56 88.44 127.72 89.56 ;
      RECT 131.04 88.44 135.64 88.6 ;
      RECT 127.56 88.44 129.36 88.6 ;
      RECT 129.08 88.36 131.27 88.52 ;
      RECT 129.08 91.4 131.27 91.56 ;
      RECT 135.48 90.36 135.64 91.48 ;
      RECT 131.04 91.32 135.64 91.48 ;
      RECT 127.56 91.32 129.36 91.48 ;
      RECT 127.56 90.36 127.72 91.48 ;
      RECT 127.56 90.36 135.64 90.52 ;
      RECT 127.56 92.8 135.64 92.96 ;
      RECT 135.48 91.84 135.64 92.96 ;
      RECT 127.56 91.84 127.72 92.96 ;
      RECT 131.04 91.84 135.64 92 ;
      RECT 127.56 91.84 129.36 92 ;
      RECT 129.08 91.76 131.27 91.92 ;
      RECT 129.08 94.8 131.27 94.96 ;
      RECT 135.48 93.76 135.64 94.88 ;
      RECT 131.04 94.72 135.64 94.88 ;
      RECT 127.56 94.72 129.36 94.88 ;
      RECT 127.56 93.76 127.72 94.88 ;
      RECT 127.56 93.76 135.64 93.92 ;
      RECT 127.56 96.2 135.64 96.36 ;
      RECT 135.48 95.24 135.64 96.36 ;
      RECT 127.56 95.24 127.72 96.36 ;
      RECT 131.04 95.24 135.64 95.4 ;
      RECT 127.56 95.24 129.36 95.4 ;
      RECT 129.08 95.16 131.27 95.32 ;
      RECT 129.08 98.2 131.27 98.36 ;
      RECT 135.48 97.16 135.64 98.28 ;
      RECT 131.04 98.12 135.64 98.28 ;
      RECT 127.56 98.12 129.36 98.28 ;
      RECT 127.56 97.16 127.72 98.28 ;
      RECT 127.56 97.16 135.64 97.32 ;
      RECT 127.56 99.6 135.64 99.76 ;
      RECT 135.48 98.64 135.64 99.76 ;
      RECT 127.56 98.64 127.72 99.76 ;
      RECT 131.04 98.64 135.64 98.8 ;
      RECT 127.56 98.64 129.36 98.8 ;
      RECT 129.08 98.56 131.27 98.72 ;
      RECT 129.08 101.6 131.27 101.76 ;
      RECT 135.48 100.56 135.64 101.68 ;
      RECT 131.04 101.52 135.64 101.68 ;
      RECT 127.56 101.52 129.36 101.68 ;
      RECT 127.56 100.56 127.72 101.68 ;
      RECT 127.56 100.56 135.64 100.72 ;
      RECT 127.56 103 135.64 103.16 ;
      RECT 135.48 102.04 135.64 103.16 ;
      RECT 127.56 102.04 127.72 103.16 ;
      RECT 131.04 102.04 135.64 102.2 ;
      RECT 127.56 102.04 129.36 102.2 ;
      RECT 129.08 101.96 131.27 102.12 ;
      RECT 129.08 105 131.27 105.16 ;
      RECT 135.48 103.96 135.64 105.08 ;
      RECT 131.04 104.92 135.64 105.08 ;
      RECT 127.56 104.92 129.36 105.08 ;
      RECT 127.56 103.96 127.72 105.08 ;
      RECT 127.56 103.96 135.64 104.12 ;
      RECT 127.56 106.4 135.64 106.56 ;
      RECT 135.48 105.44 135.64 106.56 ;
      RECT 127.56 105.44 127.72 106.56 ;
      RECT 131.04 105.44 135.64 105.6 ;
      RECT 127.56 105.44 129.36 105.6 ;
      RECT 129.08 105.36 131.27 105.52 ;
      RECT 129.08 108.4 131.27 108.56 ;
      RECT 135.48 107.36 135.64 108.48 ;
      RECT 131.04 108.32 135.64 108.48 ;
      RECT 127.56 108.32 129.36 108.48 ;
      RECT 127.56 107.36 127.72 108.48 ;
      RECT 127.56 107.36 135.64 107.52 ;
      RECT 127.56 109.8 135.64 109.96 ;
      RECT 135.48 108.84 135.64 109.96 ;
      RECT 127.56 108.84 127.72 109.96 ;
      RECT 131.04 108.84 135.64 109 ;
      RECT 127.56 108.84 129.36 109 ;
      RECT 129.08 108.76 131.27 108.92 ;
      RECT 129.08 111.8 131.27 111.96 ;
      RECT 135.48 110.76 135.64 111.88 ;
      RECT 131.04 111.72 135.64 111.88 ;
      RECT 127.56 111.72 129.36 111.88 ;
      RECT 127.56 110.76 127.72 111.88 ;
      RECT 127.56 110.76 135.64 110.92 ;
      RECT 127.56 113.2 135.64 113.36 ;
      RECT 135.48 112.24 135.64 113.36 ;
      RECT 127.56 112.24 127.72 113.36 ;
      RECT 131.04 112.24 135.64 112.4 ;
      RECT 127.56 112.24 129.36 112.4 ;
      RECT 129.08 112.16 131.27 112.32 ;
      RECT 129.08 115.2 131.27 115.36 ;
      RECT 135.48 114.16 135.64 115.28 ;
      RECT 131.04 115.12 135.64 115.28 ;
      RECT 127.56 115.12 129.36 115.28 ;
      RECT 127.56 114.16 127.72 115.28 ;
      RECT 127.56 114.16 135.64 114.32 ;
      RECT 127.56 116.6 135.64 116.76 ;
      RECT 135.48 115.64 135.64 116.76 ;
      RECT 127.56 115.64 127.72 116.76 ;
      RECT 131.04 115.64 135.64 115.8 ;
      RECT 127.56 115.64 129.36 115.8 ;
      RECT 129.08 115.56 131.27 115.72 ;
      RECT 129.08 118.6 131.27 118.76 ;
      RECT 135.48 117.56 135.64 118.68 ;
      RECT 131.04 118.52 135.64 118.68 ;
      RECT 127.56 118.52 129.36 118.68 ;
      RECT 127.56 117.56 127.72 118.68 ;
      RECT 127.56 117.56 135.64 117.72 ;
      RECT 127.56 120 135.64 120.16 ;
      RECT 135.48 119.04 135.64 120.16 ;
      RECT 127.56 119.04 127.72 120.16 ;
      RECT 131.04 119.04 135.64 119.2 ;
      RECT 127.56 119.04 129.36 119.2 ;
      RECT 129.08 118.96 131.27 119.12 ;
      RECT 129.08 122 131.27 122.16 ;
      RECT 135.48 120.96 135.64 122.08 ;
      RECT 131.04 121.92 135.64 122.08 ;
      RECT 127.56 121.92 129.36 122.08 ;
      RECT 127.56 120.96 127.72 122.08 ;
      RECT 127.56 120.96 135.64 121.12 ;
      RECT 127.56 123.4 135.64 123.56 ;
      RECT 135.48 122.44 135.64 123.56 ;
      RECT 127.56 122.44 127.72 123.56 ;
      RECT 131.04 122.44 135.64 122.6 ;
      RECT 127.56 122.44 129.36 122.6 ;
      RECT 129.08 122.36 131.27 122.52 ;
      RECT 129.08 125.4 131.27 125.56 ;
      RECT 135.48 124.36 135.64 125.48 ;
      RECT 131.04 125.32 135.64 125.48 ;
      RECT 127.56 125.32 129.36 125.48 ;
      RECT 127.56 124.36 127.72 125.48 ;
      RECT 127.56 124.36 135.64 124.52 ;
      RECT 127.56 126.8 135.64 126.96 ;
      RECT 135.48 125.84 135.64 126.96 ;
      RECT 127.56 125.84 127.72 126.96 ;
      RECT 131.04 125.84 135.64 126 ;
      RECT 127.56 125.84 129.36 126 ;
      RECT 129.08 125.76 131.27 125.92 ;
      RECT 129.08 128.8 131.27 128.96 ;
      RECT 135.48 127.76 135.64 128.88 ;
      RECT 131.04 128.72 135.64 128.88 ;
      RECT 127.56 128.72 129.36 128.88 ;
      RECT 127.56 127.76 127.72 128.88 ;
      RECT 127.56 127.76 135.64 127.92 ;
      RECT 127.56 130.2 135.64 130.36 ;
      RECT 135.48 129.24 135.64 130.36 ;
      RECT 127.56 129.24 127.72 130.36 ;
      RECT 131.04 129.24 135.64 129.4 ;
      RECT 127.56 129.24 129.36 129.4 ;
      RECT 129.08 129.16 131.27 129.32 ;
      RECT 129.08 132.2 131.27 132.36 ;
      RECT 135.48 131.16 135.64 132.28 ;
      RECT 131.04 132.12 135.64 132.28 ;
      RECT 127.56 132.12 129.36 132.28 ;
      RECT 127.56 131.16 127.72 132.28 ;
      RECT 127.56 131.16 135.64 131.32 ;
      RECT 127.56 133.6 135.64 133.76 ;
      RECT 135.48 132.64 135.64 133.76 ;
      RECT 127.56 132.64 127.72 133.76 ;
      RECT 131.04 132.64 135.64 132.8 ;
      RECT 127.56 132.64 129.36 132.8 ;
      RECT 129.08 132.56 131.27 132.72 ;
      RECT 129.08 135.6 131.27 135.76 ;
      RECT 135.48 134.56 135.64 135.68 ;
      RECT 131.04 135.52 135.64 135.68 ;
      RECT 127.56 135.52 129.36 135.68 ;
      RECT 127.56 134.56 127.72 135.68 ;
      RECT 127.56 134.56 135.64 134.72 ;
      RECT 127.56 137 135.64 137.16 ;
      RECT 135.48 136.04 135.64 137.16 ;
      RECT 127.56 136.04 127.72 137.16 ;
      RECT 131.04 136.04 135.64 136.2 ;
      RECT 127.56 136.04 129.36 136.2 ;
      RECT 129.08 135.96 131.27 136.12 ;
      RECT 129.08 139 131.27 139.16 ;
      RECT 135.48 137.96 135.64 139.08 ;
      RECT 131.04 138.92 135.64 139.08 ;
      RECT 127.56 138.92 129.36 139.08 ;
      RECT 127.56 137.96 127.72 139.08 ;
      RECT 127.56 137.96 135.64 138.12 ;
      RECT 127.56 140.4 135.64 140.56 ;
      RECT 135.48 139.44 135.64 140.56 ;
      RECT 127.56 139.44 127.72 140.56 ;
      RECT 131.04 139.44 135.64 139.6 ;
      RECT 127.56 139.44 129.36 139.6 ;
      RECT 129.08 139.36 131.27 139.52 ;
      RECT 129.08 142.4 131.27 142.56 ;
      RECT 135.48 141.36 135.64 142.48 ;
      RECT 131.04 142.32 135.64 142.48 ;
      RECT 127.56 142.32 129.36 142.48 ;
      RECT 127.56 141.36 127.72 142.48 ;
      RECT 127.56 141.36 135.64 141.52 ;
      RECT 127.56 143.8 135.64 143.96 ;
      RECT 135.48 142.84 135.64 143.96 ;
      RECT 127.56 142.84 127.72 143.96 ;
      RECT 131.04 142.84 135.64 143 ;
      RECT 127.56 142.84 129.36 143 ;
      RECT 129.08 142.76 131.27 142.92 ;
      RECT 129.08 145.8 131.27 145.96 ;
      RECT 135.48 144.76 135.64 145.88 ;
      RECT 131.04 145.72 135.64 145.88 ;
      RECT 127.56 145.72 129.36 145.88 ;
      RECT 127.56 144.76 127.72 145.88 ;
      RECT 127.56 144.76 135.64 144.92 ;
      RECT 127.56 147.2 135.64 147.36 ;
      RECT 135.48 146.24 135.64 147.36 ;
      RECT 127.56 146.24 127.72 147.36 ;
      RECT 131.04 146.24 135.64 146.4 ;
      RECT 127.56 146.24 129.36 146.4 ;
      RECT 129.08 146.16 131.27 146.32 ;
      RECT 129.08 149.2 131.27 149.36 ;
      RECT 135.48 148.16 135.64 149.28 ;
      RECT 131.04 149.12 135.64 149.28 ;
      RECT 127.56 149.12 129.36 149.28 ;
      RECT 127.56 148.16 127.72 149.28 ;
      RECT 127.56 148.16 135.64 148.32 ;
      RECT 127.56 150.6 135.64 150.76 ;
      RECT 135.48 149.64 135.64 150.76 ;
      RECT 127.56 149.64 127.72 150.76 ;
      RECT 131.04 149.64 135.64 149.8 ;
      RECT 127.56 149.64 129.36 149.8 ;
      RECT 129.08 149.56 131.27 149.72 ;
      RECT 129.08 152.6 131.27 152.76 ;
      RECT 135.48 151.56 135.64 152.68 ;
      RECT 131.04 152.52 135.64 152.68 ;
      RECT 127.56 152.52 129.36 152.68 ;
      RECT 127.56 151.56 127.72 152.68 ;
      RECT 127.56 151.56 135.64 151.72 ;
      RECT 127.56 154 135.64 154.16 ;
      RECT 135.48 153.04 135.64 154.16 ;
      RECT 127.56 153.04 127.72 154.16 ;
      RECT 131.04 153.04 135.64 153.2 ;
      RECT 127.56 153.04 129.36 153.2 ;
      RECT 129.08 152.96 131.27 153.12 ;
      RECT 129.08 156 131.27 156.16 ;
      RECT 135.48 154.96 135.64 156.08 ;
      RECT 131.04 155.92 135.64 156.08 ;
      RECT 127.56 155.92 129.36 156.08 ;
      RECT 127.56 154.96 127.72 156.08 ;
      RECT 127.56 154.96 135.64 155.12 ;
      RECT 127.56 157.4 135.64 157.56 ;
      RECT 135.48 156.44 135.64 157.56 ;
      RECT 127.56 156.44 127.72 157.56 ;
      RECT 131.04 156.44 135.64 156.6 ;
      RECT 127.56 156.44 129.36 156.6 ;
      RECT 129.08 156.36 131.27 156.52 ;
      RECT 129.08 159.4 131.27 159.56 ;
      RECT 135.48 158.36 135.64 159.48 ;
      RECT 131.04 159.32 135.64 159.48 ;
      RECT 127.56 159.32 129.36 159.48 ;
      RECT 127.56 158.36 127.72 159.48 ;
      RECT 127.56 158.36 135.64 158.52 ;
      RECT 127.56 160.8 135.64 160.96 ;
      RECT 135.48 159.84 135.64 160.96 ;
      RECT 127.56 159.84 127.72 160.96 ;
      RECT 131.04 159.84 135.64 160 ;
      RECT 127.56 159.84 129.36 160 ;
      RECT 129.08 159.76 131.27 159.92 ;
      RECT 129.08 162.8 131.27 162.96 ;
      RECT 135.48 161.76 135.64 162.88 ;
      RECT 131.04 162.72 135.64 162.88 ;
      RECT 127.56 162.72 129.36 162.88 ;
      RECT 127.56 161.76 127.72 162.88 ;
      RECT 127.56 161.76 135.64 161.92 ;
      RECT 127.56 164.2 135.64 164.36 ;
      RECT 135.48 163.24 135.64 164.36 ;
      RECT 127.56 163.24 127.72 164.36 ;
      RECT 131.04 163.24 135.64 163.4 ;
      RECT 127.56 163.24 129.36 163.4 ;
      RECT 129.08 163.16 131.27 163.32 ;
      RECT 129.08 166.2 131.27 166.36 ;
      RECT 135.48 165.16 135.64 166.28 ;
      RECT 131.04 166.12 135.64 166.28 ;
      RECT 127.56 166.12 129.36 166.28 ;
      RECT 127.56 165.16 127.72 166.28 ;
      RECT 127.56 165.16 135.64 165.32 ;
      RECT 127.56 167.6 135.64 167.76 ;
      RECT 135.48 166.64 135.64 167.76 ;
      RECT 127.56 166.64 127.72 167.76 ;
      RECT 131.04 166.64 135.64 166.8 ;
      RECT 127.56 166.64 129.36 166.8 ;
      RECT 129.08 166.56 131.27 166.72 ;
      RECT 129.08 169.6 131.27 169.76 ;
      RECT 135.48 168.56 135.64 169.68 ;
      RECT 131.04 169.52 135.64 169.68 ;
      RECT 127.56 169.52 129.36 169.68 ;
      RECT 127.56 168.56 127.72 169.68 ;
      RECT 127.56 168.56 135.64 168.72 ;
      RECT 127.56 171 135.64 171.16 ;
      RECT 135.48 170.04 135.64 171.16 ;
      RECT 127.56 170.04 127.72 171.16 ;
      RECT 131.04 170.04 135.64 170.2 ;
      RECT 127.56 170.04 129.36 170.2 ;
      RECT 129.08 169.96 131.27 170.12 ;
      RECT 129.08 173 131.27 173.16 ;
      RECT 135.48 171.96 135.64 173.08 ;
      RECT 131.04 172.92 135.64 173.08 ;
      RECT 127.56 172.92 129.36 173.08 ;
      RECT 127.56 171.96 127.72 173.08 ;
      RECT 127.56 171.96 135.64 172.12 ;
      RECT 127.56 174.4 135.64 174.56 ;
      RECT 135.48 173.44 135.64 174.56 ;
      RECT 127.56 173.44 127.72 174.56 ;
      RECT 131.04 173.44 135.64 173.6 ;
      RECT 127.56 173.44 129.36 173.6 ;
      RECT 129.08 173.36 131.27 173.52 ;
      RECT 129.08 176.4 131.27 176.56 ;
      RECT 135.48 175.36 135.64 176.48 ;
      RECT 131.04 176.32 135.64 176.48 ;
      RECT 127.56 176.32 129.36 176.48 ;
      RECT 127.56 175.36 127.72 176.48 ;
      RECT 127.56 175.36 135.64 175.52 ;
      RECT 127.56 177.8 135.64 177.96 ;
      RECT 135.48 176.84 135.64 177.96 ;
      RECT 127.56 176.84 127.72 177.96 ;
      RECT 131.04 176.84 135.64 177 ;
      RECT 127.56 176.84 129.36 177 ;
      RECT 129.08 176.76 131.27 176.92 ;
      RECT 129.08 179.8 131.27 179.96 ;
      RECT 135.48 178.76 135.64 179.88 ;
      RECT 131.04 179.72 135.64 179.88 ;
      RECT 127.56 179.72 129.36 179.88 ;
      RECT 127.56 178.76 127.72 179.88 ;
      RECT 127.56 178.76 135.64 178.92 ;
      RECT 127.56 181.2 135.64 181.36 ;
      RECT 135.48 180.24 135.64 181.36 ;
      RECT 127.56 180.24 127.72 181.36 ;
      RECT 131.04 180.24 135.64 180.4 ;
      RECT 127.56 180.24 129.36 180.4 ;
      RECT 129.08 180.16 131.27 180.32 ;
      RECT 129.08 183.2 131.27 183.36 ;
      RECT 135.48 182.16 135.64 183.28 ;
      RECT 131.04 183.12 135.64 183.28 ;
      RECT 127.56 183.12 129.36 183.28 ;
      RECT 127.56 182.16 127.72 183.28 ;
      RECT 127.56 182.16 135.64 182.32 ;
      RECT 127.56 184.6 135.64 184.76 ;
      RECT 135.48 183.64 135.64 184.76 ;
      RECT 127.56 183.64 127.72 184.76 ;
      RECT 131.04 183.64 135.64 183.8 ;
      RECT 127.56 183.64 129.36 183.8 ;
      RECT 129.08 183.56 131.27 183.72 ;
      RECT 129.08 186.6 131.27 186.76 ;
      RECT 135.48 185.56 135.64 186.68 ;
      RECT 131.04 186.52 135.64 186.68 ;
      RECT 127.56 186.52 129.36 186.68 ;
      RECT 127.56 185.56 127.72 186.68 ;
      RECT 127.56 185.56 135.64 185.72 ;
      RECT 127.56 188 135.64 188.16 ;
      RECT 135.48 187.04 135.64 188.16 ;
      RECT 127.56 187.04 127.72 188.16 ;
      RECT 131.04 187.04 135.64 187.2 ;
      RECT 127.56 187.04 129.36 187.2 ;
      RECT 129.08 186.96 131.27 187.12 ;
      RECT 129.08 190 131.27 190.16 ;
      RECT 135.48 188.96 135.64 190.08 ;
      RECT 131.04 189.92 135.64 190.08 ;
      RECT 127.56 189.92 129.36 190.08 ;
      RECT 127.56 188.96 127.72 190.08 ;
      RECT 127.56 188.96 135.64 189.12 ;
      RECT 127.56 191.4 135.64 191.56 ;
      RECT 135.48 190.44 135.64 191.56 ;
      RECT 127.56 190.44 127.72 191.56 ;
      RECT 131.04 190.44 135.64 190.6 ;
      RECT 127.56 190.44 129.36 190.6 ;
      RECT 129.08 190.36 131.27 190.52 ;
      RECT 129.08 193.4 131.27 193.56 ;
      RECT 135.48 192.36 135.64 193.48 ;
      RECT 131.04 193.32 135.64 193.48 ;
      RECT 127.56 193.32 129.36 193.48 ;
      RECT 127.56 192.36 127.72 193.48 ;
      RECT 127.56 192.36 135.64 192.52 ;
      RECT 127.56 194.8 135.64 194.96 ;
      RECT 135.48 193.84 135.64 194.96 ;
      RECT 127.56 193.84 127.72 194.96 ;
      RECT 131.04 193.84 135.64 194 ;
      RECT 127.56 193.84 129.36 194 ;
      RECT 129.08 193.76 131.27 193.92 ;
      RECT 129.08 196.8 131.27 196.96 ;
      RECT 135.48 195.76 135.64 196.88 ;
      RECT 131.04 196.72 135.64 196.88 ;
      RECT 127.56 196.72 129.36 196.88 ;
      RECT 127.56 195.76 127.72 196.88 ;
      RECT 127.56 195.76 135.64 195.92 ;
      RECT 127.56 198.2 135.64 198.36 ;
      RECT 135.48 197.24 135.64 198.36 ;
      RECT 127.56 197.24 127.72 198.36 ;
      RECT 131.04 197.24 135.64 197.4 ;
      RECT 127.56 197.24 129.36 197.4 ;
      RECT 129.08 197.16 131.27 197.32 ;
      RECT 129.08 200.2 131.27 200.36 ;
      RECT 135.48 199.16 135.64 200.28 ;
      RECT 131.04 200.12 135.64 200.28 ;
      RECT 127.56 200.12 129.36 200.28 ;
      RECT 127.56 199.16 127.72 200.28 ;
      RECT 127.56 199.16 135.64 199.32 ;
      RECT 127.56 201.6 135.64 201.76 ;
      RECT 135.48 200.64 135.64 201.76 ;
      RECT 127.56 200.64 127.72 201.76 ;
      RECT 131.04 200.64 135.64 200.8 ;
      RECT 127.56 200.64 129.36 200.8 ;
      RECT 129.08 200.56 131.27 200.72 ;
      RECT 129.08 203.6 131.27 203.76 ;
      RECT 135.48 202.56 135.64 203.68 ;
      RECT 131.04 203.52 135.64 203.68 ;
      RECT 127.56 203.52 129.36 203.68 ;
      RECT 127.56 202.56 127.72 203.68 ;
      RECT 127.56 202.56 135.64 202.72 ;
      RECT 127.56 205 135.64 205.16 ;
      RECT 135.48 204.04 135.64 205.16 ;
      RECT 127.56 204.04 127.72 205.16 ;
      RECT 131.04 204.04 135.64 204.2 ;
      RECT 127.56 204.04 129.36 204.2 ;
      RECT 129.08 203.96 131.27 204.12 ;
      RECT 129.08 207 131.27 207.16 ;
      RECT 135.48 205.96 135.64 207.08 ;
      RECT 131.04 206.92 135.64 207.08 ;
      RECT 127.56 206.92 129.36 207.08 ;
      RECT 127.56 205.96 127.72 207.08 ;
      RECT 127.56 205.96 135.64 206.12 ;
      RECT 127.56 208.4 135.64 208.56 ;
      RECT 135.48 207.44 135.64 208.56 ;
      RECT 127.56 207.44 127.72 208.56 ;
      RECT 131.04 207.44 135.64 207.6 ;
      RECT 127.56 207.44 129.36 207.6 ;
      RECT 129.08 207.36 131.27 207.52 ;
      RECT 129.08 210.4 131.27 210.56 ;
      RECT 135.48 209.36 135.64 210.48 ;
      RECT 131.04 210.32 135.64 210.48 ;
      RECT 127.56 210.32 129.36 210.48 ;
      RECT 127.56 209.36 127.72 210.48 ;
      RECT 127.56 209.36 135.64 209.52 ;
      RECT 127.56 211.8 135.64 211.96 ;
      RECT 135.48 210.84 135.64 211.96 ;
      RECT 127.56 210.84 127.72 211.96 ;
      RECT 131.04 210.84 135.64 211 ;
      RECT 127.56 210.84 129.36 211 ;
      RECT 129.08 210.76 131.27 210.92 ;
      RECT 129.08 213.8 131.27 213.96 ;
      RECT 135.48 212.76 135.64 213.88 ;
      RECT 131.04 213.72 135.64 213.88 ;
      RECT 127.56 213.72 129.36 213.88 ;
      RECT 127.56 212.76 127.72 213.88 ;
      RECT 127.56 212.76 135.64 212.92 ;
      RECT 127.56 215.2 135.64 215.36 ;
      RECT 135.48 214.24 135.64 215.36 ;
      RECT 127.56 214.24 127.72 215.36 ;
      RECT 131.04 214.24 135.64 214.4 ;
      RECT 127.56 214.24 129.36 214.4 ;
      RECT 129.08 214.16 131.27 214.32 ;
      RECT 129.08 217.2 131.27 217.36 ;
      RECT 135.48 216.16 135.64 217.28 ;
      RECT 131.04 217.12 135.64 217.28 ;
      RECT 127.56 217.12 129.36 217.28 ;
      RECT 127.56 216.16 127.72 217.28 ;
      RECT 127.56 216.16 135.64 216.32 ;
      RECT 127.56 218.6 135.64 218.76 ;
      RECT 135.48 217.64 135.64 218.76 ;
      RECT 127.56 217.64 127.72 218.76 ;
      RECT 131.04 217.64 135.64 217.8 ;
      RECT 127.56 217.64 129.36 217.8 ;
      RECT 129.08 217.56 131.27 217.72 ;
      RECT 129.08 220.6 131.27 220.76 ;
      RECT 135.48 219.56 135.64 220.68 ;
      RECT 131.04 220.52 135.64 220.68 ;
      RECT 127.56 220.52 129.36 220.68 ;
      RECT 127.56 219.56 127.72 220.68 ;
      RECT 127.56 219.56 135.64 219.72 ;
      RECT 127.56 222 135.64 222.16 ;
      RECT 135.48 221.04 135.64 222.16 ;
      RECT 127.56 221.04 127.72 222.16 ;
      RECT 131.04 221.04 135.64 221.2 ;
      RECT 127.56 221.04 129.36 221.2 ;
      RECT 129.08 220.96 131.27 221.12 ;
      RECT 129.08 224 131.27 224.16 ;
      RECT 135.48 222.96 135.64 224.08 ;
      RECT 131.04 223.92 135.64 224.08 ;
      RECT 127.56 223.92 129.36 224.08 ;
      RECT 127.56 222.96 127.72 224.08 ;
      RECT 127.56 222.96 135.64 223.12 ;
      RECT 127.56 225.4 135.64 225.56 ;
      RECT 135.48 224.44 135.64 225.56 ;
      RECT 127.56 224.44 127.72 225.56 ;
      RECT 131.04 224.44 135.64 224.6 ;
      RECT 127.56 224.44 129.36 224.6 ;
      RECT 129.08 224.36 131.27 224.52 ;
      RECT 129.08 227.4 131.27 227.56 ;
      RECT 135.48 226.36 135.64 227.48 ;
      RECT 131.04 227.32 135.64 227.48 ;
      RECT 127.56 227.32 129.36 227.48 ;
      RECT 127.56 226.36 127.72 227.48 ;
      RECT 127.56 226.36 135.64 226.52 ;
      RECT 127.56 228.8 135.64 228.96 ;
      RECT 135.48 227.84 135.64 228.96 ;
      RECT 127.56 227.84 127.72 228.96 ;
      RECT 131.04 227.84 135.64 228 ;
      RECT 127.56 227.84 129.36 228 ;
      RECT 129.08 227.76 131.27 227.92 ;
      RECT 129.08 230.8 131.27 230.96 ;
      RECT 135.48 229.76 135.64 230.88 ;
      RECT 131.04 230.72 135.64 230.88 ;
      RECT 127.56 230.72 129.36 230.88 ;
      RECT 127.56 229.76 127.72 230.88 ;
      RECT 127.56 229.76 135.64 229.92 ;
      RECT 127.56 232.2 135.64 232.36 ;
      RECT 135.48 231.24 135.64 232.36 ;
      RECT 127.56 231.24 127.72 232.36 ;
      RECT 131.04 231.24 135.64 231.4 ;
      RECT 127.56 231.24 129.36 231.4 ;
      RECT 129.08 231.16 131.27 231.32 ;
      RECT 129.08 234.2 131.27 234.36 ;
      RECT 135.48 233.16 135.64 234.28 ;
      RECT 131.04 234.12 135.64 234.28 ;
      RECT 127.56 234.12 129.36 234.28 ;
      RECT 127.56 233.16 127.72 234.28 ;
      RECT 127.56 233.16 135.64 233.32 ;
      RECT 127.56 235.6 135.64 235.76 ;
      RECT 135.48 234.64 135.64 235.76 ;
      RECT 127.56 234.64 127.72 235.76 ;
      RECT 131.04 234.64 135.64 234.8 ;
      RECT 127.56 234.64 129.36 234.8 ;
      RECT 129.08 234.56 131.27 234.72 ;
      RECT 129.08 237.6 131.27 237.76 ;
      RECT 135.48 236.56 135.64 237.68 ;
      RECT 131.04 237.52 135.64 237.68 ;
      RECT 127.56 237.52 129.36 237.68 ;
      RECT 127.56 236.56 127.72 237.68 ;
      RECT 127.56 236.56 135.64 236.72 ;
      RECT 127.56 239 135.64 239.16 ;
      RECT 135.48 238.04 135.64 239.16 ;
      RECT 127.56 238.04 127.72 239.16 ;
      RECT 131.04 238.04 135.64 238.2 ;
      RECT 127.56 238.04 129.36 238.2 ;
      RECT 129.08 237.96 131.27 238.12 ;
      RECT 129.08 241 131.27 241.16 ;
      RECT 135.48 239.96 135.64 241.08 ;
      RECT 131.04 240.92 135.64 241.08 ;
      RECT 127.56 240.92 129.36 241.08 ;
      RECT 127.56 239.96 127.72 241.08 ;
      RECT 127.56 239.96 135.64 240.12 ;
      RECT 127.56 242.4 135.64 242.56 ;
      RECT 135.48 241.44 135.64 242.56 ;
      RECT 127.56 241.44 127.72 242.56 ;
      RECT 131.04 241.44 135.64 241.6 ;
      RECT 127.56 241.44 129.36 241.6 ;
      RECT 129.08 241.36 131.27 241.52 ;
      RECT 129.08 244.4 131.27 244.56 ;
      RECT 135.48 243.36 135.64 244.48 ;
      RECT 131.04 244.32 135.64 244.48 ;
      RECT 127.56 244.32 129.36 244.48 ;
      RECT 127.56 243.36 127.72 244.48 ;
      RECT 127.56 243.36 135.64 243.52 ;
      RECT 127.56 245.8 135.64 245.96 ;
      RECT 135.48 244.84 135.64 245.96 ;
      RECT 127.56 244.84 127.72 245.96 ;
      RECT 131.04 244.84 135.64 245 ;
      RECT 127.56 244.84 129.36 245 ;
      RECT 129.08 244.76 131.27 244.92 ;
      RECT 129.08 247.8 131.27 247.96 ;
      RECT 135.48 246.76 135.64 247.88 ;
      RECT 131.04 247.72 135.64 247.88 ;
      RECT 127.56 247.72 129.36 247.88 ;
      RECT 127.56 246.76 127.72 247.88 ;
      RECT 127.56 246.76 135.64 246.92 ;
      RECT 127.56 249.2 135.64 249.36 ;
      RECT 135.48 248.24 135.64 249.36 ;
      RECT 127.56 248.24 127.72 249.36 ;
      RECT 131.04 248.24 135.64 248.4 ;
      RECT 127.56 248.24 129.36 248.4 ;
      RECT 129.08 248.16 131.27 248.32 ;
      RECT 129.08 251.2 131.27 251.36 ;
      RECT 135.48 250.16 135.64 251.28 ;
      RECT 131.04 251.12 135.64 251.28 ;
      RECT 127.56 251.12 129.36 251.28 ;
      RECT 127.56 250.16 127.72 251.28 ;
      RECT 127.56 250.16 135.64 250.32 ;
      RECT 127.56 252.6 135.64 252.76 ;
      RECT 135.48 251.64 135.64 252.76 ;
      RECT 127.56 251.64 127.72 252.76 ;
      RECT 131.04 251.64 135.64 251.8 ;
      RECT 127.56 251.64 129.36 251.8 ;
      RECT 129.08 251.56 131.27 251.72 ;
      RECT 129.08 254.6 131.27 254.76 ;
      RECT 135.48 253.56 135.64 254.68 ;
      RECT 131.04 254.52 135.64 254.68 ;
      RECT 127.56 254.52 129.36 254.68 ;
      RECT 127.56 253.56 127.72 254.68 ;
      RECT 127.56 253.56 135.64 253.72 ;
      RECT 127.56 256 135.64 256.16 ;
      RECT 135.48 255.04 135.64 256.16 ;
      RECT 127.56 255.04 127.72 256.16 ;
      RECT 131.04 255.04 135.64 255.2 ;
      RECT 127.56 255.04 129.36 255.2 ;
      RECT 129.08 254.96 131.27 255.12 ;
      RECT 129.08 258 131.27 258.16 ;
      RECT 135.48 256.96 135.64 258.08 ;
      RECT 131.04 257.92 135.64 258.08 ;
      RECT 127.56 257.92 129.36 258.08 ;
      RECT 127.56 256.96 127.72 258.08 ;
      RECT 127.56 256.96 135.64 257.12 ;
      RECT 127.56 259.4 135.64 259.56 ;
      RECT 135.48 258.44 135.64 259.56 ;
      RECT 127.56 258.44 127.72 259.56 ;
      RECT 131.04 258.44 135.64 258.6 ;
      RECT 127.56 258.44 129.36 258.6 ;
      RECT 129.08 258.36 131.27 258.52 ;
      RECT 129.08 261.4 131.27 261.56 ;
      RECT 135.48 260.36 135.64 261.48 ;
      RECT 131.04 261.32 135.64 261.48 ;
      RECT 127.56 261.32 129.36 261.48 ;
      RECT 127.56 260.36 127.72 261.48 ;
      RECT 127.56 260.36 135.64 260.52 ;
      RECT 127.56 262.8 135.64 262.96 ;
      RECT 135.48 261.84 135.64 262.96 ;
      RECT 127.56 261.84 127.72 262.96 ;
      RECT 131.04 261.84 135.64 262 ;
      RECT 127.56 261.84 129.36 262 ;
      RECT 129.08 261.76 131.27 261.92 ;
      RECT 129.08 264.8 131.27 264.96 ;
      RECT 135.48 263.76 135.64 264.88 ;
      RECT 131.04 264.72 135.64 264.88 ;
      RECT 127.56 264.72 129.36 264.88 ;
      RECT 127.56 263.76 127.72 264.88 ;
      RECT 127.56 263.76 135.64 263.92 ;
      RECT 127.56 266.2 135.64 266.36 ;
      RECT 135.48 265.24 135.64 266.36 ;
      RECT 127.56 265.24 127.72 266.36 ;
      RECT 131.04 265.24 135.64 265.4 ;
      RECT 127.56 265.24 129.36 265.4 ;
      RECT 129.08 265.16 131.27 265.32 ;
      RECT 129.08 268.2 131.27 268.36 ;
      RECT 135.48 267.16 135.64 268.28 ;
      RECT 131.04 268.12 135.64 268.28 ;
      RECT 127.56 268.12 129.36 268.28 ;
      RECT 127.56 267.16 127.72 268.28 ;
      RECT 127.56 267.16 135.64 267.32 ;
      RECT 127.56 269.6 135.64 269.76 ;
      RECT 135.48 268.64 135.64 269.76 ;
      RECT 127.56 268.64 127.72 269.76 ;
      RECT 131.04 268.64 135.64 268.8 ;
      RECT 127.56 268.64 129.36 268.8 ;
      RECT 129.08 268.56 131.27 268.72 ;
      RECT 129.08 271.6 131.27 271.76 ;
      RECT 135.48 270.56 135.64 271.68 ;
      RECT 131.04 271.52 135.64 271.68 ;
      RECT 127.56 271.52 129.36 271.68 ;
      RECT 127.56 270.56 127.72 271.68 ;
      RECT 127.56 270.56 135.64 270.72 ;
      RECT 127.56 273 135.64 273.16 ;
      RECT 135.48 272.04 135.64 273.16 ;
      RECT 127.56 272.04 127.72 273.16 ;
      RECT 131.04 272.04 135.64 272.2 ;
      RECT 127.56 272.04 129.36 272.2 ;
      RECT 129.08 271.96 131.27 272.12 ;
      RECT 129.08 275 131.27 275.16 ;
      RECT 135.48 273.96 135.64 275.08 ;
      RECT 131.04 274.92 135.64 275.08 ;
      RECT 127.56 274.92 129.36 275.08 ;
      RECT 127.56 273.96 127.72 275.08 ;
      RECT 127.56 273.96 135.64 274.12 ;
      RECT 127.56 276.4 135.64 276.56 ;
      RECT 135.48 275.44 135.64 276.56 ;
      RECT 127.56 275.44 127.72 276.56 ;
      RECT 131.04 275.44 135.64 275.6 ;
      RECT 127.56 275.44 129.36 275.6 ;
      RECT 129.08 275.36 131.27 275.52 ;
      RECT 129.08 278.4 131.27 278.56 ;
      RECT 135.48 277.36 135.64 278.48 ;
      RECT 131.04 278.32 135.64 278.48 ;
      RECT 127.56 278.32 129.36 278.48 ;
      RECT 127.56 277.36 127.72 278.48 ;
      RECT 127.56 277.36 135.64 277.52 ;
      RECT 127.56 279.8 135.64 279.96 ;
      RECT 135.48 278.84 135.64 279.96 ;
      RECT 127.56 278.84 127.72 279.96 ;
      RECT 131.04 278.84 135.64 279 ;
      RECT 127.56 278.84 129.36 279 ;
      RECT 129.08 278.76 131.27 278.92 ;
      RECT 129.08 281.8 131.27 281.96 ;
      RECT 135.48 280.76 135.64 281.88 ;
      RECT 131.04 281.72 135.64 281.88 ;
      RECT 127.56 281.72 129.36 281.88 ;
      RECT 127.56 280.76 127.72 281.88 ;
      RECT 127.56 280.76 135.64 280.92 ;
      RECT 127.56 283.2 135.64 283.36 ;
      RECT 135.48 282.24 135.64 283.36 ;
      RECT 127.56 282.24 127.72 283.36 ;
      RECT 131.04 282.24 135.64 282.4 ;
      RECT 127.56 282.24 129.36 282.4 ;
      RECT 129.08 282.16 131.27 282.32 ;
      RECT 129.08 285.2 131.27 285.36 ;
      RECT 135.48 284.16 135.64 285.28 ;
      RECT 131.04 285.12 135.64 285.28 ;
      RECT 127.56 285.12 129.36 285.28 ;
      RECT 127.56 284.16 127.72 285.28 ;
      RECT 127.56 284.16 135.64 284.32 ;
      RECT 127.56 286.6 135.64 286.76 ;
      RECT 135.48 285.64 135.64 286.76 ;
      RECT 127.56 285.64 127.72 286.76 ;
      RECT 131.04 285.64 135.64 285.8 ;
      RECT 127.56 285.64 129.36 285.8 ;
      RECT 129.08 285.56 131.27 285.72 ;
      RECT 129.08 288.6 131.27 288.76 ;
      RECT 135.48 287.56 135.64 288.68 ;
      RECT 131.04 288.52 135.64 288.68 ;
      RECT 127.56 288.52 129.36 288.68 ;
      RECT 127.56 287.56 127.72 288.68 ;
      RECT 127.56 287.56 135.64 287.72 ;
      RECT 127.56 290 135.64 290.16 ;
      RECT 135.48 289.04 135.64 290.16 ;
      RECT 127.56 289.04 127.72 290.16 ;
      RECT 131.04 289.04 135.64 289.2 ;
      RECT 127.56 289.04 129.36 289.2 ;
      RECT 129.08 288.96 131.27 289.12 ;
      RECT 129.08 292 131.27 292.16 ;
      RECT 135.48 290.96 135.64 292.08 ;
      RECT 131.04 291.92 135.64 292.08 ;
      RECT 127.56 291.92 129.36 292.08 ;
      RECT 127.56 290.96 127.72 292.08 ;
      RECT 127.56 290.96 135.64 291.12 ;
      RECT 127.56 293.4 135.64 293.56 ;
      RECT 135.48 292.44 135.64 293.56 ;
      RECT 127.56 292.44 127.72 293.56 ;
      RECT 131.04 292.44 135.64 292.6 ;
      RECT 127.56 292.44 129.36 292.6 ;
      RECT 129.08 292.36 131.27 292.52 ;
      RECT 129.08 295.4 131.27 295.56 ;
      RECT 135.48 294.36 135.64 295.48 ;
      RECT 131.04 295.32 135.64 295.48 ;
      RECT 127.56 295.32 129.36 295.48 ;
      RECT 127.56 294.36 127.72 295.48 ;
      RECT 127.56 294.36 135.64 294.52 ;
      RECT 127.56 296.8 135.64 296.96 ;
      RECT 135.48 295.84 135.64 296.96 ;
      RECT 127.56 295.84 127.72 296.96 ;
      RECT 131.04 295.84 135.64 296 ;
      RECT 127.56 295.84 129.36 296 ;
      RECT 129.08 295.76 131.27 295.92 ;
      RECT 129.08 298.8 131.27 298.96 ;
      RECT 135.48 297.76 135.64 298.88 ;
      RECT 131.04 298.72 135.64 298.88 ;
      RECT 127.56 298.72 129.36 298.88 ;
      RECT 127.56 297.76 127.72 298.88 ;
      RECT 127.56 297.76 135.64 297.92 ;
      RECT 127.56 300.2 135.64 300.36 ;
      RECT 135.48 299.24 135.64 300.36 ;
      RECT 127.56 299.24 127.72 300.36 ;
      RECT 131.04 299.24 135.64 299.4 ;
      RECT 127.56 299.24 129.36 299.4 ;
      RECT 129.08 299.16 131.27 299.32 ;
      RECT 129.08 302.2 131.27 302.36 ;
      RECT 135.48 301.16 135.64 302.28 ;
      RECT 131.04 302.12 135.64 302.28 ;
      RECT 127.56 302.12 129.36 302.28 ;
      RECT 127.56 301.16 127.72 302.28 ;
      RECT 127.56 301.16 135.64 301.32 ;
      RECT 127.56 303.6 135.64 303.76 ;
      RECT 135.48 302.64 135.64 303.76 ;
      RECT 127.56 302.64 127.72 303.76 ;
      RECT 131.04 302.64 135.64 302.8 ;
      RECT 127.56 302.64 129.36 302.8 ;
      RECT 129.08 302.56 131.27 302.72 ;
      RECT 129.08 305.6 131.27 305.76 ;
      RECT 135.48 304.56 135.64 305.68 ;
      RECT 131.04 305.52 135.64 305.68 ;
      RECT 127.56 305.52 129.36 305.68 ;
      RECT 127.56 304.56 127.72 305.68 ;
      RECT 127.56 304.56 135.64 304.72 ;
      RECT 127.56 307 135.64 307.16 ;
      RECT 135.48 306.04 135.64 307.16 ;
      RECT 127.56 306.04 127.72 307.16 ;
      RECT 131.04 306.04 135.64 306.2 ;
      RECT 127.56 306.04 129.36 306.2 ;
      RECT 129.08 305.96 131.27 306.12 ;
      RECT 129.08 309 131.27 309.16 ;
      RECT 135.48 307.96 135.64 309.08 ;
      RECT 131.04 308.92 135.64 309.08 ;
      RECT 127.56 308.92 129.36 309.08 ;
      RECT 127.56 307.96 127.72 309.08 ;
      RECT 127.56 307.96 135.64 308.12 ;
      RECT 127.56 310.4 135.64 310.56 ;
      RECT 135.48 309.44 135.64 310.56 ;
      RECT 127.56 309.44 127.72 310.56 ;
      RECT 131.04 309.44 135.64 309.6 ;
      RECT 127.56 309.44 129.36 309.6 ;
      RECT 129.08 309.36 131.27 309.52 ;
      RECT 129.08 312.4 131.27 312.56 ;
      RECT 135.48 311.36 135.64 312.48 ;
      RECT 131.04 312.32 135.64 312.48 ;
      RECT 127.56 312.32 129.36 312.48 ;
      RECT 127.56 311.36 127.72 312.48 ;
      RECT 127.56 311.36 135.64 311.52 ;
      RECT 127.56 313.8 135.64 313.96 ;
      RECT 135.48 312.84 135.64 313.96 ;
      RECT 127.56 312.84 127.72 313.96 ;
      RECT 131.04 312.84 135.64 313 ;
      RECT 127.56 312.84 129.36 313 ;
      RECT 129.08 312.76 131.27 312.92 ;
      RECT 129.08 315.8 131.27 315.96 ;
      RECT 135.48 314.76 135.64 315.88 ;
      RECT 131.04 315.72 135.64 315.88 ;
      RECT 127.56 315.72 129.36 315.88 ;
      RECT 127.56 314.76 127.72 315.88 ;
      RECT 127.56 314.76 135.64 314.92 ;
      RECT 127.56 317.2 135.64 317.36 ;
      RECT 135.48 316.24 135.64 317.36 ;
      RECT 127.56 316.24 127.72 317.36 ;
      RECT 131.04 316.24 135.64 316.4 ;
      RECT 127.56 316.24 129.36 316.4 ;
      RECT 129.08 316.16 131.27 316.32 ;
      RECT 129.08 319.2 131.27 319.36 ;
      RECT 135.48 318.16 135.64 319.28 ;
      RECT 131.04 319.12 135.64 319.28 ;
      RECT 127.56 319.12 129.36 319.28 ;
      RECT 127.56 318.16 127.72 319.28 ;
      RECT 127.56 318.16 135.64 318.32 ;
      RECT 127.56 320.6 135.64 320.76 ;
      RECT 135.48 319.64 135.64 320.76 ;
      RECT 127.56 319.64 127.72 320.76 ;
      RECT 131.04 319.64 135.64 319.8 ;
      RECT 127.56 319.64 129.36 319.8 ;
      RECT 129.08 319.56 131.27 319.72 ;
      RECT 129.08 322.6 131.27 322.76 ;
      RECT 135.48 321.56 135.64 322.68 ;
      RECT 131.04 322.52 135.64 322.68 ;
      RECT 127.56 322.52 129.36 322.68 ;
      RECT 127.56 321.56 127.72 322.68 ;
      RECT 127.56 321.56 135.64 321.72 ;
      RECT 127.56 324 135.64 324.16 ;
      RECT 135.48 323.04 135.64 324.16 ;
      RECT 127.56 323.04 127.72 324.16 ;
      RECT 131.04 323.04 135.64 323.2 ;
      RECT 127.56 323.04 129.36 323.2 ;
      RECT 129.08 322.96 131.27 323.12 ;
      RECT 129.08 326 131.27 326.16 ;
      RECT 135.48 324.96 135.64 326.08 ;
      RECT 131.04 325.92 135.64 326.08 ;
      RECT 127.56 325.92 129.36 326.08 ;
      RECT 127.56 324.96 127.72 326.08 ;
      RECT 127.56 324.96 135.64 325.12 ;
      RECT 127.56 327.4 135.64 327.56 ;
      RECT 135.48 326.44 135.64 327.56 ;
      RECT 127.56 326.44 127.72 327.56 ;
      RECT 131.04 326.44 135.64 326.6 ;
      RECT 127.56 326.44 129.36 326.6 ;
      RECT 129.08 326.36 131.27 326.52 ;
      RECT 129.08 329.4 131.27 329.56 ;
      RECT 135.48 328.36 135.64 329.48 ;
      RECT 131.04 329.32 135.64 329.48 ;
      RECT 127.56 329.32 129.36 329.48 ;
      RECT 127.56 328.36 127.72 329.48 ;
      RECT 127.56 328.36 135.64 328.52 ;
      RECT 127.56 330.8 135.64 330.96 ;
      RECT 135.48 329.84 135.64 330.96 ;
      RECT 127.56 329.84 127.72 330.96 ;
      RECT 131.04 329.84 135.64 330 ;
      RECT 127.56 329.84 129.36 330 ;
      RECT 129.08 329.76 131.27 329.92 ;
      RECT 129.08 332.8 131.27 332.96 ;
      RECT 135.48 331.76 135.64 332.88 ;
      RECT 131.04 332.72 135.64 332.88 ;
      RECT 127.56 332.72 129.36 332.88 ;
      RECT 127.56 331.76 127.72 332.88 ;
      RECT 127.56 331.76 135.64 331.92 ;
      RECT 127.56 334.2 135.64 334.36 ;
      RECT 135.48 333.24 135.64 334.36 ;
      RECT 127.56 333.24 127.72 334.36 ;
      RECT 131.04 333.24 135.64 333.4 ;
      RECT 127.56 333.24 129.36 333.4 ;
      RECT 129.08 333.16 131.27 333.32 ;
      RECT 129.08 336.2 131.27 336.36 ;
      RECT 135.48 335.16 135.64 336.28 ;
      RECT 131.04 336.12 135.64 336.28 ;
      RECT 127.56 336.12 129.36 336.28 ;
      RECT 127.56 335.16 127.72 336.28 ;
      RECT 127.56 335.16 135.64 335.32 ;
      RECT 127.56 337.6 135.64 337.76 ;
      RECT 135.48 336.64 135.64 337.76 ;
      RECT 127.56 336.64 127.72 337.76 ;
      RECT 131.04 336.64 135.64 336.8 ;
      RECT 127.56 336.64 129.36 336.8 ;
      RECT 129.08 336.56 131.27 336.72 ;
      RECT 129.08 339.6 131.27 339.76 ;
      RECT 135.48 338.56 135.64 339.68 ;
      RECT 131.04 339.52 135.64 339.68 ;
      RECT 127.56 339.52 129.36 339.68 ;
      RECT 127.56 338.56 127.72 339.68 ;
      RECT 127.56 338.56 135.64 338.72 ;
      RECT 127.56 341 135.64 341.16 ;
      RECT 135.48 340.04 135.64 341.16 ;
      RECT 127.56 340.04 127.72 341.16 ;
      RECT 131.04 340.04 135.64 340.2 ;
      RECT 127.56 340.04 129.36 340.2 ;
      RECT 129.08 339.96 131.27 340.12 ;
      RECT 129.08 343 131.27 343.16 ;
      RECT 135.48 341.96 135.64 343.08 ;
      RECT 131.04 342.92 135.64 343.08 ;
      RECT 127.56 342.92 129.36 343.08 ;
      RECT 127.56 341.96 127.72 343.08 ;
      RECT 127.56 341.96 135.64 342.12 ;
      RECT 127.56 344.4 135.64 344.56 ;
      RECT 135.48 343.44 135.64 344.56 ;
      RECT 127.56 343.44 127.72 344.56 ;
      RECT 131.04 343.44 135.64 343.6 ;
      RECT 127.56 343.44 129.36 343.6 ;
      RECT 129.08 343.36 131.27 343.52 ;
      RECT 129.08 346.4 131.27 346.56 ;
      RECT 135.48 345.36 135.64 346.48 ;
      RECT 131.04 346.32 135.64 346.48 ;
      RECT 127.56 346.32 129.36 346.48 ;
      RECT 127.56 345.36 127.72 346.48 ;
      RECT 127.56 345.36 135.64 345.52 ;
      RECT 127.56 347.8 135.64 347.96 ;
      RECT 135.48 346.84 135.64 347.96 ;
      RECT 127.56 346.84 127.72 347.96 ;
      RECT 131.04 346.84 135.64 347 ;
      RECT 127.56 346.84 129.36 347 ;
      RECT 129.08 346.76 131.27 346.92 ;
      RECT 129.08 349.8 131.27 349.96 ;
      RECT 135.48 348.76 135.64 349.88 ;
      RECT 131.04 349.72 135.64 349.88 ;
      RECT 127.56 349.72 129.36 349.88 ;
      RECT 127.56 348.76 127.72 349.88 ;
      RECT 127.56 348.76 135.64 348.92 ;
      RECT 127.56 351.2 135.64 351.36 ;
      RECT 135.48 350.24 135.64 351.36 ;
      RECT 127.56 350.24 127.72 351.36 ;
      RECT 131.04 350.24 135.64 350.4 ;
      RECT 127.56 350.24 129.36 350.4 ;
      RECT 129.08 350.16 131.27 350.32 ;
      RECT 129.08 353.2 131.27 353.36 ;
      RECT 135.48 352.16 135.64 353.28 ;
      RECT 131.04 353.12 135.64 353.28 ;
      RECT 127.56 353.12 129.36 353.28 ;
      RECT 127.56 352.16 127.72 353.28 ;
      RECT 127.56 352.16 135.64 352.32 ;
      RECT 127.56 354.6 135.64 354.76 ;
      RECT 135.48 353.64 135.64 354.76 ;
      RECT 127.56 353.64 127.72 354.76 ;
      RECT 131.04 353.64 135.64 353.8 ;
      RECT 127.56 353.64 129.36 353.8 ;
      RECT 129.08 353.56 131.27 353.72 ;
      RECT 129.08 356.6 131.27 356.76 ;
      RECT 135.48 355.56 135.64 356.68 ;
      RECT 131.04 356.52 135.64 356.68 ;
      RECT 127.56 356.52 129.36 356.68 ;
      RECT 127.56 355.56 127.72 356.68 ;
      RECT 127.56 355.56 135.64 355.72 ;
      RECT 127.56 358 135.64 358.16 ;
      RECT 135.48 357.04 135.64 358.16 ;
      RECT 127.56 357.04 127.72 358.16 ;
      RECT 131.04 357.04 135.64 357.2 ;
      RECT 127.56 357.04 129.36 357.2 ;
      RECT 129.08 356.96 131.27 357.12 ;
      RECT 129.08 360 131.27 360.16 ;
      RECT 135.48 358.96 135.64 360.08 ;
      RECT 131.04 359.92 135.64 360.08 ;
      RECT 127.56 359.92 129.36 360.08 ;
      RECT 127.56 358.96 127.72 360.08 ;
      RECT 127.56 358.96 135.64 359.12 ;
      RECT 127.56 361.4 135.64 361.56 ;
      RECT 135.48 360.44 135.64 361.56 ;
      RECT 127.56 360.44 127.72 361.56 ;
      RECT 131.04 360.44 135.64 360.6 ;
      RECT 127.56 360.44 129.36 360.6 ;
      RECT 129.08 360.36 131.27 360.52 ;
      RECT 129.08 363.4 131.27 363.56 ;
      RECT 135.48 362.36 135.64 363.48 ;
      RECT 131.04 363.32 135.64 363.48 ;
      RECT 127.56 363.32 129.36 363.48 ;
      RECT 127.56 362.36 127.72 363.48 ;
      RECT 127.56 362.36 135.64 362.52 ;
      RECT 127.56 364.8 135.64 364.96 ;
      RECT 135.48 363.84 135.64 364.96 ;
      RECT 127.56 363.84 127.72 364.96 ;
      RECT 131.04 363.84 135.64 364 ;
      RECT 127.56 363.84 129.36 364 ;
      RECT 129.08 363.76 131.27 363.92 ;
      RECT 129.08 366.8 131.27 366.96 ;
      RECT 135.48 365.76 135.64 366.88 ;
      RECT 131.04 366.72 135.64 366.88 ;
      RECT 127.56 366.72 129.36 366.88 ;
      RECT 127.56 365.76 127.72 366.88 ;
      RECT 127.56 365.76 135.64 365.92 ;
      RECT 127.56 368.2 135.64 368.36 ;
      RECT 135.48 367.24 135.64 368.36 ;
      RECT 127.56 367.24 127.72 368.36 ;
      RECT 131.04 367.24 135.64 367.4 ;
      RECT 127.56 367.24 129.36 367.4 ;
      RECT 129.08 367.16 131.27 367.32 ;
      RECT 129.08 370.2 131.27 370.36 ;
      RECT 135.48 369.16 135.64 370.28 ;
      RECT 131.04 370.12 135.64 370.28 ;
      RECT 127.56 370.12 129.36 370.28 ;
      RECT 127.56 369.16 127.72 370.28 ;
      RECT 127.56 369.16 135.64 369.32 ;
      RECT 127.56 371.6 135.64 371.76 ;
      RECT 135.48 370.64 135.64 371.76 ;
      RECT 127.56 370.64 127.72 371.76 ;
      RECT 131.04 370.64 135.64 370.8 ;
      RECT 127.56 370.64 129.36 370.8 ;
      RECT 129.08 370.56 131.27 370.72 ;
      RECT 129.08 373.6 131.27 373.76 ;
      RECT 135.48 372.56 135.64 373.68 ;
      RECT 131.04 373.52 135.64 373.68 ;
      RECT 127.56 373.52 129.36 373.68 ;
      RECT 127.56 372.56 127.72 373.68 ;
      RECT 127.56 372.56 135.64 372.72 ;
      RECT 127.56 375 135.64 375.16 ;
      RECT 135.48 374.04 135.64 375.16 ;
      RECT 127.56 374.04 127.72 375.16 ;
      RECT 131.04 374.04 135.64 374.2 ;
      RECT 127.56 374.04 129.36 374.2 ;
      RECT 129.08 373.96 131.27 374.12 ;
      RECT 129.08 377 131.27 377.16 ;
      RECT 135.48 375.96 135.64 377.08 ;
      RECT 131.04 376.92 135.64 377.08 ;
      RECT 127.56 376.92 129.36 377.08 ;
      RECT 127.56 375.96 127.72 377.08 ;
      RECT 127.56 375.96 135.64 376.12 ;
      RECT 127.56 378.4 135.64 378.56 ;
      RECT 135.48 377.44 135.64 378.56 ;
      RECT 127.56 377.44 127.72 378.56 ;
      RECT 131.04 377.44 135.64 377.6 ;
      RECT 127.56 377.44 129.36 377.6 ;
      RECT 129.08 377.36 131.27 377.52 ;
      RECT 129.08 380.4 131.27 380.56 ;
      RECT 135.48 379.36 135.64 380.48 ;
      RECT 131.04 380.32 135.64 380.48 ;
      RECT 127.56 380.32 129.36 380.48 ;
      RECT 127.56 379.36 127.72 380.48 ;
      RECT 127.56 379.36 135.64 379.52 ;
      RECT 127.56 381.8 135.64 381.96 ;
      RECT 135.48 380.84 135.64 381.96 ;
      RECT 127.56 380.84 127.72 381.96 ;
      RECT 131.04 380.84 135.64 381 ;
      RECT 127.56 380.84 129.36 381 ;
      RECT 129.08 380.76 131.27 380.92 ;
      RECT 129.08 383.8 131.27 383.96 ;
      RECT 135.48 382.76 135.64 383.88 ;
      RECT 131.04 383.72 135.64 383.88 ;
      RECT 127.56 383.72 129.36 383.88 ;
      RECT 127.56 382.76 127.72 383.88 ;
      RECT 127.56 382.76 135.64 382.92 ;
      RECT 127.56 385.2 135.64 385.36 ;
      RECT 135.48 384.24 135.64 385.36 ;
      RECT 127.56 384.24 127.72 385.36 ;
      RECT 131.04 384.24 135.64 384.4 ;
      RECT 127.56 384.24 129.36 384.4 ;
      RECT 129.08 384.16 131.27 384.32 ;
      RECT 129.08 387.2 131.27 387.36 ;
      RECT 135.48 386.16 135.64 387.28 ;
      RECT 131.04 387.12 135.64 387.28 ;
      RECT 127.56 387.12 129.36 387.28 ;
      RECT 127.56 386.16 127.72 387.28 ;
      RECT 127.56 386.16 135.64 386.32 ;
      RECT 127.56 388.6 135.64 388.76 ;
      RECT 135.48 387.64 135.64 388.76 ;
      RECT 127.56 387.64 127.72 388.76 ;
      RECT 131.04 387.64 135.64 387.8 ;
      RECT 127.56 387.64 129.36 387.8 ;
      RECT 129.08 387.56 131.27 387.72 ;
      RECT 129.08 390.6 131.27 390.76 ;
      RECT 135.48 389.56 135.64 390.68 ;
      RECT 131.04 390.52 135.64 390.68 ;
      RECT 127.56 390.52 129.36 390.68 ;
      RECT 127.56 389.56 127.72 390.68 ;
      RECT 127.56 389.56 135.64 389.72 ;
      RECT 127.56 392 135.64 392.16 ;
      RECT 135.48 391.04 135.64 392.16 ;
      RECT 127.56 391.04 127.72 392.16 ;
      RECT 131.04 391.04 135.64 391.2 ;
      RECT 127.56 391.04 129.36 391.2 ;
      RECT 129.08 390.96 131.27 391.12 ;
      RECT 129.08 394 131.27 394.16 ;
      RECT 135.48 392.96 135.64 394.08 ;
      RECT 131.04 393.92 135.64 394.08 ;
      RECT 127.56 393.92 129.36 394.08 ;
      RECT 127.56 392.96 127.72 394.08 ;
      RECT 127.56 392.96 135.64 393.12 ;
      RECT 127.56 395.4 135.64 395.56 ;
      RECT 135.48 394.44 135.64 395.56 ;
      RECT 127.56 394.44 127.72 395.56 ;
      RECT 131.04 394.44 135.64 394.6 ;
      RECT 127.56 394.44 129.36 394.6 ;
      RECT 129.08 394.36 131.27 394.52 ;
      RECT 129.08 397.4 131.27 397.56 ;
      RECT 135.48 396.36 135.64 397.48 ;
      RECT 131.04 397.32 135.64 397.48 ;
      RECT 127.56 397.32 129.36 397.48 ;
      RECT 127.56 396.36 127.72 397.48 ;
      RECT 127.56 396.36 135.64 396.52 ;
      RECT 127.56 398.8 135.64 398.96 ;
      RECT 135.48 397.84 135.64 398.96 ;
      RECT 127.56 397.84 127.72 398.96 ;
      RECT 131.04 397.84 135.64 398 ;
      RECT 127.56 397.84 129.36 398 ;
      RECT 129.08 397.76 131.27 397.92 ;
      RECT 129.08 400.8 131.27 400.96 ;
      RECT 135.48 399.76 135.64 400.88 ;
      RECT 131.04 400.72 135.64 400.88 ;
      RECT 127.56 400.72 129.36 400.88 ;
      RECT 127.56 399.76 127.72 400.88 ;
      RECT 127.56 399.76 135.64 399.92 ;
      RECT 127.56 402.2 135.64 402.36 ;
      RECT 135.48 401.24 135.64 402.36 ;
      RECT 127.56 401.24 127.72 402.36 ;
      RECT 131.04 401.24 135.64 401.4 ;
      RECT 127.56 401.24 129.36 401.4 ;
      RECT 129.08 401.16 131.27 401.32 ;
      RECT 129.08 404.2 131.27 404.36 ;
      RECT 135.48 403.16 135.64 404.28 ;
      RECT 131.04 404.12 135.64 404.28 ;
      RECT 127.56 404.12 129.36 404.28 ;
      RECT 127.56 403.16 127.72 404.28 ;
      RECT 127.56 403.16 135.64 403.32 ;
      RECT 127.56 405.6 135.64 405.76 ;
      RECT 135.48 404.64 135.64 405.76 ;
      RECT 127.56 404.64 127.72 405.76 ;
      RECT 131.04 404.64 135.64 404.8 ;
      RECT 127.56 404.64 129.36 404.8 ;
      RECT 129.08 404.56 131.27 404.72 ;
      RECT 129.08 407.6 131.27 407.76 ;
      RECT 135.48 406.56 135.64 407.68 ;
      RECT 131.04 407.52 135.64 407.68 ;
      RECT 127.56 407.52 129.36 407.68 ;
      RECT 127.56 406.56 127.72 407.68 ;
      RECT 127.56 406.56 135.64 406.72 ;
      RECT 127.56 409 135.64 409.16 ;
      RECT 135.48 408.04 135.64 409.16 ;
      RECT 127.56 408.04 127.72 409.16 ;
      RECT 131.04 408.04 135.64 408.2 ;
      RECT 127.56 408.04 129.36 408.2 ;
      RECT 129.08 407.96 131.27 408.12 ;
      RECT 129.08 411 131.27 411.16 ;
      RECT 135.48 409.96 135.64 411.08 ;
      RECT 131.04 410.92 135.64 411.08 ;
      RECT 127.56 410.92 129.36 411.08 ;
      RECT 127.56 409.96 127.72 411.08 ;
      RECT 127.56 409.96 135.64 410.12 ;
      RECT 127.56 412.4 135.64 412.56 ;
      RECT 135.48 411.44 135.64 412.56 ;
      RECT 127.56 411.44 127.72 412.56 ;
      RECT 131.04 411.44 135.64 411.6 ;
      RECT 127.56 411.44 129.36 411.6 ;
      RECT 129.08 411.36 131.27 411.52 ;
      RECT 129.08 414.4 131.27 414.56 ;
      RECT 135.48 413.36 135.64 414.48 ;
      RECT 131.04 414.32 135.64 414.48 ;
      RECT 127.56 414.32 129.36 414.48 ;
      RECT 127.56 413.36 127.72 414.48 ;
      RECT 127.56 413.36 135.64 413.52 ;
      RECT 127.56 415.8 135.64 415.96 ;
      RECT 135.48 414.84 135.64 415.96 ;
      RECT 127.56 414.84 127.72 415.96 ;
      RECT 131.04 414.84 135.64 415 ;
      RECT 127.56 414.84 129.36 415 ;
      RECT 129.08 414.76 131.27 414.92 ;
      RECT 129.08 417.8 131.27 417.96 ;
      RECT 135.48 416.76 135.64 417.88 ;
      RECT 131.04 417.72 135.64 417.88 ;
      RECT 127.56 417.72 129.36 417.88 ;
      RECT 127.56 416.76 127.72 417.88 ;
      RECT 127.56 416.76 135.64 416.92 ;
      RECT 127.56 419.2 135.64 419.36 ;
      RECT 135.48 418.24 135.64 419.36 ;
      RECT 127.56 418.24 127.72 419.36 ;
      RECT 131.04 418.24 135.64 418.4 ;
      RECT 127.56 418.24 129.36 418.4 ;
      RECT 129.08 418.16 131.27 418.32 ;
      RECT 129.08 421.2 131.27 421.36 ;
      RECT 135.48 420.16 135.64 421.28 ;
      RECT 131.04 421.12 135.64 421.28 ;
      RECT 127.56 421.12 129.36 421.28 ;
      RECT 127.56 420.16 127.72 421.28 ;
      RECT 127.56 420.16 135.64 420.32 ;
      RECT 127.56 422.6 135.64 422.76 ;
      RECT 135.48 421.64 135.64 422.76 ;
      RECT 127.56 421.64 127.72 422.76 ;
      RECT 131.04 421.64 135.64 421.8 ;
      RECT 127.56 421.64 129.36 421.8 ;
      RECT 129.08 421.56 131.27 421.72 ;
      RECT 129.08 424.6 131.27 424.76 ;
      RECT 135.48 423.56 135.64 424.68 ;
      RECT 131.04 424.52 135.64 424.68 ;
      RECT 127.56 424.52 129.36 424.68 ;
      RECT 127.56 423.56 127.72 424.68 ;
      RECT 127.56 423.56 135.64 423.72 ;
      RECT 127.56 426 135.64 426.16 ;
      RECT 135.48 425.04 135.64 426.16 ;
      RECT 127.56 425.04 127.72 426.16 ;
      RECT 131.04 425.04 135.64 425.2 ;
      RECT 127.56 425.04 129.36 425.2 ;
      RECT 129.08 424.96 131.27 425.12 ;
      RECT 129.08 428 131.27 428.16 ;
      RECT 135.48 426.96 135.64 428.08 ;
      RECT 131.04 427.92 135.64 428.08 ;
      RECT 127.56 427.92 129.36 428.08 ;
      RECT 127.56 426.96 127.72 428.08 ;
      RECT 127.56 426.96 135.64 427.12 ;
      RECT 127.56 429.4 135.64 429.56 ;
      RECT 135.48 428.44 135.64 429.56 ;
      RECT 127.56 428.44 127.72 429.56 ;
      RECT 131.04 428.44 135.64 428.6 ;
      RECT 127.56 428.44 129.36 428.6 ;
      RECT 129.08 428.36 131.27 428.52 ;
      RECT 129.08 431.4 131.27 431.56 ;
      RECT 135.48 430.36 135.64 431.48 ;
      RECT 131.04 431.32 135.64 431.48 ;
      RECT 127.56 431.32 129.36 431.48 ;
      RECT 127.56 430.36 127.72 431.48 ;
      RECT 127.56 430.36 135.64 430.52 ;
      RECT 127.56 432.8 135.64 432.96 ;
      RECT 135.48 431.84 135.64 432.96 ;
      RECT 127.56 431.84 127.72 432.96 ;
      RECT 131.04 431.84 135.64 432 ;
      RECT 127.56 431.84 129.36 432 ;
      RECT 129.08 431.76 131.27 431.92 ;
      RECT 129.08 434.8 131.27 434.96 ;
      RECT 135.48 433.76 135.64 434.88 ;
      RECT 131.04 434.72 135.64 434.88 ;
      RECT 127.56 434.72 129.36 434.88 ;
      RECT 127.56 433.76 127.72 434.88 ;
      RECT 127.56 433.76 135.64 433.92 ;
      RECT 127.56 436.2 135.64 436.36 ;
      RECT 135.48 435.24 135.64 436.36 ;
      RECT 127.56 435.24 127.72 436.36 ;
      RECT 131.04 435.24 135.64 435.4 ;
      RECT 127.56 435.24 129.36 435.4 ;
      RECT 129.08 435.16 131.27 435.32 ;
      RECT 129.08 438.2 131.27 438.36 ;
      RECT 135.48 437.16 135.64 438.28 ;
      RECT 131.04 438.12 135.64 438.28 ;
      RECT 127.56 438.12 129.36 438.28 ;
      RECT 127.56 437.16 127.72 438.28 ;
      RECT 127.56 437.16 135.64 437.32 ;
      RECT 127.56 439.6 135.64 439.76 ;
      RECT 135.48 438.64 135.64 439.76 ;
      RECT 127.56 438.64 127.72 439.76 ;
      RECT 131.04 438.64 135.64 438.8 ;
      RECT 127.56 438.64 129.36 438.8 ;
      RECT 129.08 438.56 131.27 438.72 ;
      RECT 129.08 441.6 131.27 441.76 ;
      RECT 135.48 440.56 135.64 441.68 ;
      RECT 131.04 441.52 135.64 441.68 ;
      RECT 127.56 441.52 129.36 441.68 ;
      RECT 127.56 440.56 127.72 441.68 ;
      RECT 127.56 440.56 135.64 440.72 ;
      RECT 127.56 443 135.64 443.16 ;
      RECT 135.48 442.04 135.64 443.16 ;
      RECT 127.56 442.04 127.72 443.16 ;
      RECT 131.04 442.04 135.64 442.2 ;
      RECT 127.56 442.04 129.36 442.2 ;
      RECT 129.08 441.96 131.27 442.12 ;
      RECT 129.08 445 131.27 445.16 ;
      RECT 135.48 443.96 135.64 445.08 ;
      RECT 131.04 444.92 135.64 445.08 ;
      RECT 127.56 444.92 129.36 445.08 ;
      RECT 127.56 443.96 127.72 445.08 ;
      RECT 127.56 443.96 135.64 444.12 ;
      RECT 127.56 446.4 135.64 446.56 ;
      RECT 135.48 445.44 135.64 446.56 ;
      RECT 127.56 445.44 127.72 446.56 ;
      RECT 131.04 445.44 135.64 445.6 ;
      RECT 127.56 445.44 129.36 445.6 ;
      RECT 129.08 445.36 131.27 445.52 ;
      RECT 129.08 448.4 131.27 448.56 ;
      RECT 135.48 447.36 135.64 448.48 ;
      RECT 131.04 448.32 135.64 448.48 ;
      RECT 127.56 448.32 129.36 448.48 ;
      RECT 127.56 447.36 127.72 448.48 ;
      RECT 127.56 447.36 135.64 447.52 ;
      RECT 127.56 449.8 135.64 449.96 ;
      RECT 135.48 448.84 135.64 449.96 ;
      RECT 127.56 448.84 127.72 449.96 ;
      RECT 131.04 448.84 135.64 449 ;
      RECT 127.56 448.84 129.36 449 ;
      RECT 129.08 448.76 131.27 448.92 ;
      RECT 129.08 451.8 131.27 451.96 ;
      RECT 135.48 450.76 135.64 451.88 ;
      RECT 131.04 451.72 135.64 451.88 ;
      RECT 127.56 451.72 129.36 451.88 ;
      RECT 127.56 450.76 127.72 451.88 ;
      RECT 127.56 450.76 135.64 450.92 ;
      RECT 127.56 453.2 135.64 453.36 ;
      RECT 135.48 452.24 135.64 453.36 ;
      RECT 127.56 452.24 127.72 453.36 ;
      RECT 131.04 452.24 135.64 452.4 ;
      RECT 127.56 452.24 129.36 452.4 ;
      RECT 129.08 452.16 131.27 452.32 ;
      RECT 129.08 455.2 131.27 455.36 ;
      RECT 135.48 454.16 135.64 455.28 ;
      RECT 131.04 455.12 135.64 455.28 ;
      RECT 127.56 455.12 129.36 455.28 ;
      RECT 127.56 454.16 127.72 455.28 ;
      RECT 127.56 454.16 135.64 454.32 ;
      RECT 127.56 456.6 135.64 456.76 ;
      RECT 135.48 455.64 135.64 456.76 ;
      RECT 127.56 455.64 127.72 456.76 ;
      RECT 131.04 455.64 135.64 455.8 ;
      RECT 127.56 455.64 129.36 455.8 ;
      RECT 129.08 455.56 131.27 455.72 ;
      RECT 129.08 458.6 131.27 458.76 ;
      RECT 135.48 457.56 135.64 458.68 ;
      RECT 131.04 458.52 135.64 458.68 ;
      RECT 127.56 458.52 129.36 458.68 ;
      RECT 127.56 457.56 127.72 458.68 ;
      RECT 127.56 457.56 135.64 457.72 ;
      RECT 127.56 460 135.64 460.16 ;
      RECT 135.48 459.04 135.64 460.16 ;
      RECT 127.56 459.04 127.72 460.16 ;
      RECT 131.04 459.04 135.64 459.2 ;
      RECT 127.56 459.04 129.36 459.2 ;
      RECT 129.08 458.96 131.27 459.12 ;
      RECT 129.08 462 131.27 462.16 ;
      RECT 135.48 460.96 135.64 462.08 ;
      RECT 131.04 461.92 135.64 462.08 ;
      RECT 127.56 461.92 129.36 462.08 ;
      RECT 127.56 460.96 127.72 462.08 ;
      RECT 127.56 460.96 135.64 461.12 ;
      RECT 127.56 463.4 135.64 463.56 ;
      RECT 135.48 462.44 135.64 463.56 ;
      RECT 127.56 462.44 127.72 463.56 ;
      RECT 131.04 462.44 135.64 462.6 ;
      RECT 127.56 462.44 129.36 462.6 ;
      RECT 129.08 462.36 131.27 462.52 ;
      RECT 129.08 465.4 131.27 465.56 ;
      RECT 135.48 464.36 135.64 465.48 ;
      RECT 131.04 465.32 135.64 465.48 ;
      RECT 127.56 465.32 129.36 465.48 ;
      RECT 127.56 464.36 127.72 465.48 ;
      RECT 127.56 464.36 135.64 464.52 ;
      RECT 127.56 466.8 135.64 466.96 ;
      RECT 135.48 465.84 135.64 466.96 ;
      RECT 127.56 465.84 127.72 466.96 ;
      RECT 131.04 465.84 135.64 466 ;
      RECT 127.56 465.84 129.36 466 ;
      RECT 129.08 465.76 131.27 465.92 ;
      RECT 129.08 468.8 131.27 468.96 ;
      RECT 135.48 467.76 135.64 468.88 ;
      RECT 131.04 468.72 135.64 468.88 ;
      RECT 127.56 468.72 129.36 468.88 ;
      RECT 127.56 467.76 127.72 468.88 ;
      RECT 127.56 467.76 135.64 467.92 ;
      RECT 127.56 470.2 135.64 470.36 ;
      RECT 135.48 469.24 135.64 470.36 ;
      RECT 127.56 469.24 127.72 470.36 ;
      RECT 131.04 469.24 135.64 469.4 ;
      RECT 127.56 469.24 129.36 469.4 ;
      RECT 129.08 469.16 131.27 469.32 ;
      RECT 129.08 472.2 131.27 472.36 ;
      RECT 135.48 471.16 135.64 472.28 ;
      RECT 131.04 472.12 135.64 472.28 ;
      RECT 127.56 472.12 129.36 472.28 ;
      RECT 127.56 471.16 127.72 472.28 ;
      RECT 127.56 471.16 135.64 471.32 ;
      RECT 127.56 473.6 135.64 473.76 ;
      RECT 135.48 472.64 135.64 473.76 ;
      RECT 127.56 472.64 127.72 473.76 ;
      RECT 131.04 472.64 135.64 472.8 ;
      RECT 127.56 472.64 129.36 472.8 ;
      RECT 129.08 472.56 131.27 472.72 ;
      RECT 129.08 475.6 131.27 475.76 ;
      RECT 135.48 474.56 135.64 475.68 ;
      RECT 131.04 475.52 135.64 475.68 ;
      RECT 127.56 475.52 129.36 475.68 ;
      RECT 127.56 474.56 127.72 475.68 ;
      RECT 127.56 474.56 135.64 474.72 ;
      RECT 127.56 477 135.64 477.16 ;
      RECT 135.48 476.04 135.64 477.16 ;
      RECT 127.56 476.04 127.72 477.16 ;
      RECT 131.04 476.04 135.64 476.2 ;
      RECT 127.56 476.04 129.36 476.2 ;
      RECT 129.08 475.96 131.27 476.12 ;
      RECT 129.08 479 131.27 479.16 ;
      RECT 135.48 477.96 135.64 479.08 ;
      RECT 131.04 478.92 135.64 479.08 ;
      RECT 127.56 478.92 129.36 479.08 ;
      RECT 127.56 477.96 127.72 479.08 ;
      RECT 127.56 477.96 135.64 478.12 ;
      RECT 127.56 480.4 135.64 480.56 ;
      RECT 135.48 479.44 135.64 480.56 ;
      RECT 127.56 479.44 127.72 480.56 ;
      RECT 131.04 479.44 135.64 479.6 ;
      RECT 127.56 479.44 129.36 479.6 ;
      RECT 129.08 479.36 131.27 479.52 ;
      RECT 129.08 482.4 131.27 482.56 ;
      RECT 135.48 481.36 135.64 482.48 ;
      RECT 131.04 482.32 135.64 482.48 ;
      RECT 127.56 482.32 129.36 482.48 ;
      RECT 127.56 481.36 127.72 482.48 ;
      RECT 127.56 481.36 135.64 481.52 ;
      RECT 127.56 483.8 135.64 483.96 ;
      RECT 135.48 482.84 135.64 483.96 ;
      RECT 127.56 482.84 127.72 483.96 ;
      RECT 131.04 482.84 135.64 483 ;
      RECT 127.56 482.84 129.36 483 ;
      RECT 129.08 482.76 131.27 482.92 ;
      RECT 129.08 485.8 131.27 485.96 ;
      RECT 135.48 484.76 135.64 485.88 ;
      RECT 131.04 485.72 135.64 485.88 ;
      RECT 127.56 485.72 129.36 485.88 ;
      RECT 127.56 484.76 127.72 485.88 ;
      RECT 127.56 484.76 135.64 484.92 ;
      RECT 127.56 487.2 135.64 487.36 ;
      RECT 135.48 486.24 135.64 487.36 ;
      RECT 127.56 486.24 127.72 487.36 ;
      RECT 131.04 486.24 135.64 486.4 ;
      RECT 127.56 486.24 129.36 486.4 ;
      RECT 129.08 486.16 131.27 486.32 ;
      RECT 129.08 489.2 131.27 489.36 ;
      RECT 135.48 488.16 135.64 489.28 ;
      RECT 131.04 489.12 135.64 489.28 ;
      RECT 127.56 489.12 129.36 489.28 ;
      RECT 127.56 488.16 127.72 489.28 ;
      RECT 127.56 488.16 135.64 488.32 ;
      RECT 127.56 490.6 135.64 490.76 ;
      RECT 135.48 489.64 135.64 490.76 ;
      RECT 127.56 489.64 127.72 490.76 ;
      RECT 131.04 489.64 135.64 489.8 ;
      RECT 127.56 489.64 129.36 489.8 ;
      RECT 129.08 489.56 131.27 489.72 ;
      RECT 129.08 492.6 131.27 492.76 ;
      RECT 135.48 491.56 135.64 492.68 ;
      RECT 131.04 492.52 135.64 492.68 ;
      RECT 127.56 492.52 129.36 492.68 ;
      RECT 127.56 491.56 127.72 492.68 ;
      RECT 127.56 491.56 135.64 491.72 ;
      RECT 127.56 494 135.64 494.16 ;
      RECT 135.48 493.04 135.64 494.16 ;
      RECT 127.56 493.04 127.72 494.16 ;
      RECT 131.04 493.04 135.64 493.2 ;
      RECT 127.56 493.04 129.36 493.2 ;
      RECT 129.08 492.96 131.27 493.12 ;
      RECT 129.08 496 131.27 496.16 ;
      RECT 135.48 494.96 135.64 496.08 ;
      RECT 131.04 495.92 135.64 496.08 ;
      RECT 127.56 495.92 129.36 496.08 ;
      RECT 127.56 494.96 127.72 496.08 ;
      RECT 127.56 494.96 135.64 495.12 ;
      RECT 127.56 497.4 135.64 497.56 ;
      RECT 135.48 496.44 135.64 497.56 ;
      RECT 127.56 496.44 127.72 497.56 ;
      RECT 131.04 496.44 135.64 496.6 ;
      RECT 127.56 496.44 129.36 496.6 ;
      RECT 129.08 496.36 131.27 496.52 ;
      RECT 129.08 499.4 131.27 499.56 ;
      RECT 135.48 498.36 135.64 499.48 ;
      RECT 131.04 499.32 135.64 499.48 ;
      RECT 127.56 499.32 129.36 499.48 ;
      RECT 127.56 498.36 127.72 499.48 ;
      RECT 127.56 498.36 135.64 498.52 ;
      RECT 127.56 500.8 135.64 500.96 ;
      RECT 135.48 499.84 135.64 500.96 ;
      RECT 127.56 499.84 127.72 500.96 ;
      RECT 131.04 499.84 135.64 500 ;
      RECT 127.56 499.84 129.36 500 ;
      RECT 129.08 499.76 131.27 499.92 ;
      RECT 129.08 502.8 131.27 502.96 ;
      RECT 135.48 501.76 135.64 502.88 ;
      RECT 131.04 502.72 135.64 502.88 ;
      RECT 127.56 502.72 129.36 502.88 ;
      RECT 127.56 501.76 127.72 502.88 ;
      RECT 127.56 501.76 135.64 501.92 ;
      RECT 127.56 504.2 135.64 504.36 ;
      RECT 135.48 503.24 135.64 504.36 ;
      RECT 127.56 503.24 127.72 504.36 ;
      RECT 131.04 503.24 135.64 503.4 ;
      RECT 127.56 503.24 129.36 503.4 ;
      RECT 129.08 503.16 131.27 503.32 ;
      RECT 135.11 14.52 135.27 16.86 ;
      RECT 135.24 13.22 135.4 14.84 ;
      RECT 135.11 31.09 135.27 35.75 ;
      RECT 135.11 32.25 135.37 32.53 ;
      RECT 133.33 26.46 135.35 26.62 ;
      RECT 133.33 25.35 133.49 26.62 ;
      RECT 133.41 22.91 133.57 25.51 ;
      RECT 133.41 56.46 133.57 59.14 ;
      RECT 133.33 55.49 133.49 56.62 ;
      RECT 133.33 55.49 135.35 55.65 ;
      RECT 135.11 49.75 135.31 51.3 ;
      RECT 135.11 46.54 135.27 51.3 ;
      RECT 133.99 55.09 135.25 55.25 ;
      RECT 133.99 49.77 134.15 55.25 ;
      RECT 133.27 49.77 134.15 49.93 ;
      RECT 133.27 32.48 133.43 49.93 ;
      RECT 133.27 45.9 134.09 46.06 ;
      RECT 133.27 36.23 134.09 36.39 ;
      RECT 133.27 32.48 134.15 32.64 ;
      RECT 133.99 27.04 134.15 32.64 ;
      RECT 133.99 27.04 135.25 27.2 ;
      RECT 134.37 45.9 135.17 46.06 ;
      RECT 135.01 44.89 135.17 46.06 ;
      RECT 135.03 38.57 135.19 45.17 ;
      RECT 134.23 38.57 134.39 45.17 ;
      RECT 134.23 38.57 134.69 38.73 ;
      RECT 134.53 36.23 134.69 38.73 ;
      RECT 134.37 36.23 135.05 36.39 ;
      RECT 130.74 70.44 130.96 70.72 ;
      RECT 130.74 70.44 134.79 70.6 ;
      RECT 130.74 71.92 134.79 72.08 ;
      RECT 130.74 71.8 130.96 72.08 ;
      RECT 130.74 73.84 130.96 74.12 ;
      RECT 130.74 73.84 134.79 74 ;
      RECT 130.74 75.32 134.79 75.48 ;
      RECT 130.74 75.2 130.96 75.48 ;
      RECT 130.74 77.24 130.96 77.52 ;
      RECT 130.74 77.24 134.79 77.4 ;
      RECT 130.74 78.72 134.79 78.88 ;
      RECT 130.74 78.6 130.96 78.88 ;
      RECT 130.74 80.64 130.96 80.92 ;
      RECT 130.74 80.64 134.79 80.8 ;
      RECT 130.74 82.12 134.79 82.28 ;
      RECT 130.74 82 130.96 82.28 ;
      RECT 130.74 84.04 130.96 84.32 ;
      RECT 130.74 84.04 134.79 84.2 ;
      RECT 130.74 85.52 134.79 85.68 ;
      RECT 130.74 85.4 130.96 85.68 ;
      RECT 130.74 87.44 130.96 87.72 ;
      RECT 130.74 87.44 134.79 87.6 ;
      RECT 130.74 88.92 134.79 89.08 ;
      RECT 130.74 88.8 130.96 89.08 ;
      RECT 130.74 90.84 130.96 91.12 ;
      RECT 130.74 90.84 134.79 91 ;
      RECT 130.74 92.32 134.79 92.48 ;
      RECT 130.74 92.2 130.96 92.48 ;
      RECT 130.74 94.24 130.96 94.52 ;
      RECT 130.74 94.24 134.79 94.4 ;
      RECT 130.74 95.72 134.79 95.88 ;
      RECT 130.74 95.6 130.96 95.88 ;
      RECT 130.74 97.64 130.96 97.92 ;
      RECT 130.74 97.64 134.79 97.8 ;
      RECT 130.74 99.12 134.79 99.28 ;
      RECT 130.74 99 130.96 99.28 ;
      RECT 130.74 101.04 130.96 101.32 ;
      RECT 130.74 101.04 134.79 101.2 ;
      RECT 130.74 102.52 134.79 102.68 ;
      RECT 130.74 102.4 130.96 102.68 ;
      RECT 130.74 104.44 130.96 104.72 ;
      RECT 130.74 104.44 134.79 104.6 ;
      RECT 130.74 105.92 134.79 106.08 ;
      RECT 130.74 105.8 130.96 106.08 ;
      RECT 130.74 107.84 130.96 108.12 ;
      RECT 130.74 107.84 134.79 108 ;
      RECT 130.74 109.32 134.79 109.48 ;
      RECT 130.74 109.2 130.96 109.48 ;
      RECT 130.74 111.24 130.96 111.52 ;
      RECT 130.74 111.24 134.79 111.4 ;
      RECT 130.74 112.72 134.79 112.88 ;
      RECT 130.74 112.6 130.96 112.88 ;
      RECT 130.74 114.64 130.96 114.92 ;
      RECT 130.74 114.64 134.79 114.8 ;
      RECT 130.74 116.12 134.79 116.28 ;
      RECT 130.74 116 130.96 116.28 ;
      RECT 130.74 118.04 130.96 118.32 ;
      RECT 130.74 118.04 134.79 118.2 ;
      RECT 130.74 119.52 134.79 119.68 ;
      RECT 130.74 119.4 130.96 119.68 ;
      RECT 130.74 121.44 130.96 121.72 ;
      RECT 130.74 121.44 134.79 121.6 ;
      RECT 130.74 122.92 134.79 123.08 ;
      RECT 130.74 122.8 130.96 123.08 ;
      RECT 130.74 124.84 130.96 125.12 ;
      RECT 130.74 124.84 134.79 125 ;
      RECT 130.74 126.32 134.79 126.48 ;
      RECT 130.74 126.2 130.96 126.48 ;
      RECT 130.74 128.24 130.96 128.52 ;
      RECT 130.74 128.24 134.79 128.4 ;
      RECT 130.74 129.72 134.79 129.88 ;
      RECT 130.74 129.6 130.96 129.88 ;
      RECT 130.74 131.64 130.96 131.92 ;
      RECT 130.74 131.64 134.79 131.8 ;
      RECT 130.74 133.12 134.79 133.28 ;
      RECT 130.74 133 130.96 133.28 ;
      RECT 130.74 135.04 130.96 135.32 ;
      RECT 130.74 135.04 134.79 135.2 ;
      RECT 130.74 136.52 134.79 136.68 ;
      RECT 130.74 136.4 130.96 136.68 ;
      RECT 130.74 138.44 130.96 138.72 ;
      RECT 130.74 138.44 134.79 138.6 ;
      RECT 130.74 139.92 134.79 140.08 ;
      RECT 130.74 139.8 130.96 140.08 ;
      RECT 130.74 141.84 130.96 142.12 ;
      RECT 130.74 141.84 134.79 142 ;
      RECT 130.74 143.32 134.79 143.48 ;
      RECT 130.74 143.2 130.96 143.48 ;
      RECT 130.74 145.24 130.96 145.52 ;
      RECT 130.74 145.24 134.79 145.4 ;
      RECT 130.74 146.72 134.79 146.88 ;
      RECT 130.74 146.6 130.96 146.88 ;
      RECT 130.74 148.64 130.96 148.92 ;
      RECT 130.74 148.64 134.79 148.8 ;
      RECT 130.74 150.12 134.79 150.28 ;
      RECT 130.74 150 130.96 150.28 ;
      RECT 130.74 152.04 130.96 152.32 ;
      RECT 130.74 152.04 134.79 152.2 ;
      RECT 130.74 153.52 134.79 153.68 ;
      RECT 130.74 153.4 130.96 153.68 ;
      RECT 130.74 155.44 130.96 155.72 ;
      RECT 130.74 155.44 134.79 155.6 ;
      RECT 130.74 156.92 134.79 157.08 ;
      RECT 130.74 156.8 130.96 157.08 ;
      RECT 130.74 158.84 130.96 159.12 ;
      RECT 130.74 158.84 134.79 159 ;
      RECT 130.74 160.32 134.79 160.48 ;
      RECT 130.74 160.2 130.96 160.48 ;
      RECT 130.74 162.24 130.96 162.52 ;
      RECT 130.74 162.24 134.79 162.4 ;
      RECT 130.74 163.72 134.79 163.88 ;
      RECT 130.74 163.6 130.96 163.88 ;
      RECT 130.74 165.64 130.96 165.92 ;
      RECT 130.74 165.64 134.79 165.8 ;
      RECT 130.74 167.12 134.79 167.28 ;
      RECT 130.74 167 130.96 167.28 ;
      RECT 130.74 169.04 130.96 169.32 ;
      RECT 130.74 169.04 134.79 169.2 ;
      RECT 130.74 170.52 134.79 170.68 ;
      RECT 130.74 170.4 130.96 170.68 ;
      RECT 130.74 172.44 130.96 172.72 ;
      RECT 130.74 172.44 134.79 172.6 ;
      RECT 130.74 173.92 134.79 174.08 ;
      RECT 130.74 173.8 130.96 174.08 ;
      RECT 130.74 175.84 130.96 176.12 ;
      RECT 130.74 175.84 134.79 176 ;
      RECT 130.74 177.32 134.79 177.48 ;
      RECT 130.74 177.2 130.96 177.48 ;
      RECT 130.74 179.24 130.96 179.52 ;
      RECT 130.74 179.24 134.79 179.4 ;
      RECT 130.74 180.72 134.79 180.88 ;
      RECT 130.74 180.6 130.96 180.88 ;
      RECT 130.74 182.64 130.96 182.92 ;
      RECT 130.74 182.64 134.79 182.8 ;
      RECT 130.74 184.12 134.79 184.28 ;
      RECT 130.74 184 130.96 184.28 ;
      RECT 130.74 186.04 130.96 186.32 ;
      RECT 130.74 186.04 134.79 186.2 ;
      RECT 130.74 187.52 134.79 187.68 ;
      RECT 130.74 187.4 130.96 187.68 ;
      RECT 130.74 189.44 130.96 189.72 ;
      RECT 130.74 189.44 134.79 189.6 ;
      RECT 130.74 190.92 134.79 191.08 ;
      RECT 130.74 190.8 130.96 191.08 ;
      RECT 130.74 192.84 130.96 193.12 ;
      RECT 130.74 192.84 134.79 193 ;
      RECT 130.74 194.32 134.79 194.48 ;
      RECT 130.74 194.2 130.96 194.48 ;
      RECT 130.74 196.24 130.96 196.52 ;
      RECT 130.74 196.24 134.79 196.4 ;
      RECT 130.74 197.72 134.79 197.88 ;
      RECT 130.74 197.6 130.96 197.88 ;
      RECT 130.74 199.64 130.96 199.92 ;
      RECT 130.74 199.64 134.79 199.8 ;
      RECT 130.74 201.12 134.79 201.28 ;
      RECT 130.74 201 130.96 201.28 ;
      RECT 130.74 203.04 130.96 203.32 ;
      RECT 130.74 203.04 134.79 203.2 ;
      RECT 130.74 204.52 134.79 204.68 ;
      RECT 130.74 204.4 130.96 204.68 ;
      RECT 130.74 206.44 130.96 206.72 ;
      RECT 130.74 206.44 134.79 206.6 ;
      RECT 130.74 207.92 134.79 208.08 ;
      RECT 130.74 207.8 130.96 208.08 ;
      RECT 130.74 209.84 130.96 210.12 ;
      RECT 130.74 209.84 134.79 210 ;
      RECT 130.74 211.32 134.79 211.48 ;
      RECT 130.74 211.2 130.96 211.48 ;
      RECT 130.74 213.24 130.96 213.52 ;
      RECT 130.74 213.24 134.79 213.4 ;
      RECT 130.74 214.72 134.79 214.88 ;
      RECT 130.74 214.6 130.96 214.88 ;
      RECT 130.74 216.64 130.96 216.92 ;
      RECT 130.74 216.64 134.79 216.8 ;
      RECT 130.74 218.12 134.79 218.28 ;
      RECT 130.74 218 130.96 218.28 ;
      RECT 130.74 220.04 130.96 220.32 ;
      RECT 130.74 220.04 134.79 220.2 ;
      RECT 130.74 221.52 134.79 221.68 ;
      RECT 130.74 221.4 130.96 221.68 ;
      RECT 130.74 223.44 130.96 223.72 ;
      RECT 130.74 223.44 134.79 223.6 ;
      RECT 130.74 224.92 134.79 225.08 ;
      RECT 130.74 224.8 130.96 225.08 ;
      RECT 130.74 226.84 130.96 227.12 ;
      RECT 130.74 226.84 134.79 227 ;
      RECT 130.74 228.32 134.79 228.48 ;
      RECT 130.74 228.2 130.96 228.48 ;
      RECT 130.74 230.24 130.96 230.52 ;
      RECT 130.74 230.24 134.79 230.4 ;
      RECT 130.74 231.72 134.79 231.88 ;
      RECT 130.74 231.6 130.96 231.88 ;
      RECT 130.74 233.64 130.96 233.92 ;
      RECT 130.74 233.64 134.79 233.8 ;
      RECT 130.74 235.12 134.79 235.28 ;
      RECT 130.74 235 130.96 235.28 ;
      RECT 130.74 237.04 130.96 237.32 ;
      RECT 130.74 237.04 134.79 237.2 ;
      RECT 130.74 238.52 134.79 238.68 ;
      RECT 130.74 238.4 130.96 238.68 ;
      RECT 130.74 240.44 130.96 240.72 ;
      RECT 130.74 240.44 134.79 240.6 ;
      RECT 130.74 241.92 134.79 242.08 ;
      RECT 130.74 241.8 130.96 242.08 ;
      RECT 130.74 243.84 130.96 244.12 ;
      RECT 130.74 243.84 134.79 244 ;
      RECT 130.74 245.32 134.79 245.48 ;
      RECT 130.74 245.2 130.96 245.48 ;
      RECT 130.74 247.24 130.96 247.52 ;
      RECT 130.74 247.24 134.79 247.4 ;
      RECT 130.74 248.72 134.79 248.88 ;
      RECT 130.74 248.6 130.96 248.88 ;
      RECT 130.74 250.64 130.96 250.92 ;
      RECT 130.74 250.64 134.79 250.8 ;
      RECT 130.74 252.12 134.79 252.28 ;
      RECT 130.74 252 130.96 252.28 ;
      RECT 130.74 254.04 130.96 254.32 ;
      RECT 130.74 254.04 134.79 254.2 ;
      RECT 130.74 255.52 134.79 255.68 ;
      RECT 130.74 255.4 130.96 255.68 ;
      RECT 130.74 257.44 130.96 257.72 ;
      RECT 130.74 257.44 134.79 257.6 ;
      RECT 130.74 258.92 134.79 259.08 ;
      RECT 130.74 258.8 130.96 259.08 ;
      RECT 130.74 260.84 130.96 261.12 ;
      RECT 130.74 260.84 134.79 261 ;
      RECT 130.74 262.32 134.79 262.48 ;
      RECT 130.74 262.2 130.96 262.48 ;
      RECT 130.74 264.24 130.96 264.52 ;
      RECT 130.74 264.24 134.79 264.4 ;
      RECT 130.74 265.72 134.79 265.88 ;
      RECT 130.74 265.6 130.96 265.88 ;
      RECT 130.74 267.64 130.96 267.92 ;
      RECT 130.74 267.64 134.79 267.8 ;
      RECT 130.74 269.12 134.79 269.28 ;
      RECT 130.74 269 130.96 269.28 ;
      RECT 130.74 271.04 130.96 271.32 ;
      RECT 130.74 271.04 134.79 271.2 ;
      RECT 130.74 272.52 134.79 272.68 ;
      RECT 130.74 272.4 130.96 272.68 ;
      RECT 130.74 274.44 130.96 274.72 ;
      RECT 130.74 274.44 134.79 274.6 ;
      RECT 130.74 275.92 134.79 276.08 ;
      RECT 130.74 275.8 130.96 276.08 ;
      RECT 130.74 277.84 130.96 278.12 ;
      RECT 130.74 277.84 134.79 278 ;
      RECT 130.74 279.32 134.79 279.48 ;
      RECT 130.74 279.2 130.96 279.48 ;
      RECT 130.74 281.24 130.96 281.52 ;
      RECT 130.74 281.24 134.79 281.4 ;
      RECT 130.74 282.72 134.79 282.88 ;
      RECT 130.74 282.6 130.96 282.88 ;
      RECT 130.74 284.64 130.96 284.92 ;
      RECT 130.74 284.64 134.79 284.8 ;
      RECT 130.74 286.12 134.79 286.28 ;
      RECT 130.74 286 130.96 286.28 ;
      RECT 130.74 288.04 130.96 288.32 ;
      RECT 130.74 288.04 134.79 288.2 ;
      RECT 130.74 289.52 134.79 289.68 ;
      RECT 130.74 289.4 130.96 289.68 ;
      RECT 130.74 291.44 130.96 291.72 ;
      RECT 130.74 291.44 134.79 291.6 ;
      RECT 130.74 292.92 134.79 293.08 ;
      RECT 130.74 292.8 130.96 293.08 ;
      RECT 130.74 294.84 130.96 295.12 ;
      RECT 130.74 294.84 134.79 295 ;
      RECT 130.74 296.32 134.79 296.48 ;
      RECT 130.74 296.2 130.96 296.48 ;
      RECT 130.74 298.24 130.96 298.52 ;
      RECT 130.74 298.24 134.79 298.4 ;
      RECT 130.74 299.72 134.79 299.88 ;
      RECT 130.74 299.6 130.96 299.88 ;
      RECT 130.74 301.64 130.96 301.92 ;
      RECT 130.74 301.64 134.79 301.8 ;
      RECT 130.74 303.12 134.79 303.28 ;
      RECT 130.74 303 130.96 303.28 ;
      RECT 130.74 305.04 130.96 305.32 ;
      RECT 130.74 305.04 134.79 305.2 ;
      RECT 130.74 306.52 134.79 306.68 ;
      RECT 130.74 306.4 130.96 306.68 ;
      RECT 130.74 308.44 130.96 308.72 ;
      RECT 130.74 308.44 134.79 308.6 ;
      RECT 130.74 309.92 134.79 310.08 ;
      RECT 130.74 309.8 130.96 310.08 ;
      RECT 130.74 311.84 130.96 312.12 ;
      RECT 130.74 311.84 134.79 312 ;
      RECT 130.74 313.32 134.79 313.48 ;
      RECT 130.74 313.2 130.96 313.48 ;
      RECT 130.74 315.24 130.96 315.52 ;
      RECT 130.74 315.24 134.79 315.4 ;
      RECT 130.74 316.72 134.79 316.88 ;
      RECT 130.74 316.6 130.96 316.88 ;
      RECT 130.74 318.64 130.96 318.92 ;
      RECT 130.74 318.64 134.79 318.8 ;
      RECT 130.74 320.12 134.79 320.28 ;
      RECT 130.74 320 130.96 320.28 ;
      RECT 130.74 322.04 130.96 322.32 ;
      RECT 130.74 322.04 134.79 322.2 ;
      RECT 130.74 323.52 134.79 323.68 ;
      RECT 130.74 323.4 130.96 323.68 ;
      RECT 130.74 325.44 130.96 325.72 ;
      RECT 130.74 325.44 134.79 325.6 ;
      RECT 130.74 326.92 134.79 327.08 ;
      RECT 130.74 326.8 130.96 327.08 ;
      RECT 130.74 328.84 130.96 329.12 ;
      RECT 130.74 328.84 134.79 329 ;
      RECT 130.74 330.32 134.79 330.48 ;
      RECT 130.74 330.2 130.96 330.48 ;
      RECT 130.74 332.24 130.96 332.52 ;
      RECT 130.74 332.24 134.79 332.4 ;
      RECT 130.74 333.72 134.79 333.88 ;
      RECT 130.74 333.6 130.96 333.88 ;
      RECT 130.74 335.64 130.96 335.92 ;
      RECT 130.74 335.64 134.79 335.8 ;
      RECT 130.74 337.12 134.79 337.28 ;
      RECT 130.74 337 130.96 337.28 ;
      RECT 130.74 339.04 130.96 339.32 ;
      RECT 130.74 339.04 134.79 339.2 ;
      RECT 130.74 340.52 134.79 340.68 ;
      RECT 130.74 340.4 130.96 340.68 ;
      RECT 130.74 342.44 130.96 342.72 ;
      RECT 130.74 342.44 134.79 342.6 ;
      RECT 130.74 343.92 134.79 344.08 ;
      RECT 130.74 343.8 130.96 344.08 ;
      RECT 130.74 345.84 130.96 346.12 ;
      RECT 130.74 345.84 134.79 346 ;
      RECT 130.74 347.32 134.79 347.48 ;
      RECT 130.74 347.2 130.96 347.48 ;
      RECT 130.74 349.24 130.96 349.52 ;
      RECT 130.74 349.24 134.79 349.4 ;
      RECT 130.74 350.72 134.79 350.88 ;
      RECT 130.74 350.6 130.96 350.88 ;
      RECT 130.74 352.64 130.96 352.92 ;
      RECT 130.74 352.64 134.79 352.8 ;
      RECT 130.74 354.12 134.79 354.28 ;
      RECT 130.74 354 130.96 354.28 ;
      RECT 130.74 356.04 130.96 356.32 ;
      RECT 130.74 356.04 134.79 356.2 ;
      RECT 130.74 357.52 134.79 357.68 ;
      RECT 130.74 357.4 130.96 357.68 ;
      RECT 130.74 359.44 130.96 359.72 ;
      RECT 130.74 359.44 134.79 359.6 ;
      RECT 130.74 360.92 134.79 361.08 ;
      RECT 130.74 360.8 130.96 361.08 ;
      RECT 130.74 362.84 130.96 363.12 ;
      RECT 130.74 362.84 134.79 363 ;
      RECT 130.74 364.32 134.79 364.48 ;
      RECT 130.74 364.2 130.96 364.48 ;
      RECT 130.74 366.24 130.96 366.52 ;
      RECT 130.74 366.24 134.79 366.4 ;
      RECT 130.74 367.72 134.79 367.88 ;
      RECT 130.74 367.6 130.96 367.88 ;
      RECT 130.74 369.64 130.96 369.92 ;
      RECT 130.74 369.64 134.79 369.8 ;
      RECT 130.74 371.12 134.79 371.28 ;
      RECT 130.74 371 130.96 371.28 ;
      RECT 130.74 373.04 130.96 373.32 ;
      RECT 130.74 373.04 134.79 373.2 ;
      RECT 130.74 374.52 134.79 374.68 ;
      RECT 130.74 374.4 130.96 374.68 ;
      RECT 130.74 376.44 130.96 376.72 ;
      RECT 130.74 376.44 134.79 376.6 ;
      RECT 130.74 377.92 134.79 378.08 ;
      RECT 130.74 377.8 130.96 378.08 ;
      RECT 130.74 379.84 130.96 380.12 ;
      RECT 130.74 379.84 134.79 380 ;
      RECT 130.74 381.32 134.79 381.48 ;
      RECT 130.74 381.2 130.96 381.48 ;
      RECT 130.74 383.24 130.96 383.52 ;
      RECT 130.74 383.24 134.79 383.4 ;
      RECT 130.74 384.72 134.79 384.88 ;
      RECT 130.74 384.6 130.96 384.88 ;
      RECT 130.74 386.64 130.96 386.92 ;
      RECT 130.74 386.64 134.79 386.8 ;
      RECT 130.74 388.12 134.79 388.28 ;
      RECT 130.74 388 130.96 388.28 ;
      RECT 130.74 390.04 130.96 390.32 ;
      RECT 130.74 390.04 134.79 390.2 ;
      RECT 130.74 391.52 134.79 391.68 ;
      RECT 130.74 391.4 130.96 391.68 ;
      RECT 130.74 393.44 130.96 393.72 ;
      RECT 130.74 393.44 134.79 393.6 ;
      RECT 130.74 394.92 134.79 395.08 ;
      RECT 130.74 394.8 130.96 395.08 ;
      RECT 130.74 396.84 130.96 397.12 ;
      RECT 130.74 396.84 134.79 397 ;
      RECT 130.74 398.32 134.79 398.48 ;
      RECT 130.74 398.2 130.96 398.48 ;
      RECT 130.74 400.24 130.96 400.52 ;
      RECT 130.74 400.24 134.79 400.4 ;
      RECT 130.74 401.72 134.79 401.88 ;
      RECT 130.74 401.6 130.96 401.88 ;
      RECT 130.74 403.64 130.96 403.92 ;
      RECT 130.74 403.64 134.79 403.8 ;
      RECT 130.74 405.12 134.79 405.28 ;
      RECT 130.74 405 130.96 405.28 ;
      RECT 130.74 407.04 130.96 407.32 ;
      RECT 130.74 407.04 134.79 407.2 ;
      RECT 130.74 408.52 134.79 408.68 ;
      RECT 130.74 408.4 130.96 408.68 ;
      RECT 130.74 410.44 130.96 410.72 ;
      RECT 130.74 410.44 134.79 410.6 ;
      RECT 130.74 411.92 134.79 412.08 ;
      RECT 130.74 411.8 130.96 412.08 ;
      RECT 130.74 413.84 130.96 414.12 ;
      RECT 130.74 413.84 134.79 414 ;
      RECT 130.74 415.32 134.79 415.48 ;
      RECT 130.74 415.2 130.96 415.48 ;
      RECT 130.74 417.24 130.96 417.52 ;
      RECT 130.74 417.24 134.79 417.4 ;
      RECT 130.74 418.72 134.79 418.88 ;
      RECT 130.74 418.6 130.96 418.88 ;
      RECT 130.74 420.64 130.96 420.92 ;
      RECT 130.74 420.64 134.79 420.8 ;
      RECT 130.74 422.12 134.79 422.28 ;
      RECT 130.74 422 130.96 422.28 ;
      RECT 130.74 424.04 130.96 424.32 ;
      RECT 130.74 424.04 134.79 424.2 ;
      RECT 130.74 425.52 134.79 425.68 ;
      RECT 130.74 425.4 130.96 425.68 ;
      RECT 130.74 427.44 130.96 427.72 ;
      RECT 130.74 427.44 134.79 427.6 ;
      RECT 130.74 428.92 134.79 429.08 ;
      RECT 130.74 428.8 130.96 429.08 ;
      RECT 130.74 430.84 130.96 431.12 ;
      RECT 130.74 430.84 134.79 431 ;
      RECT 130.74 432.32 134.79 432.48 ;
      RECT 130.74 432.2 130.96 432.48 ;
      RECT 130.74 434.24 130.96 434.52 ;
      RECT 130.74 434.24 134.79 434.4 ;
      RECT 130.74 435.72 134.79 435.88 ;
      RECT 130.74 435.6 130.96 435.88 ;
      RECT 130.74 437.64 130.96 437.92 ;
      RECT 130.74 437.64 134.79 437.8 ;
      RECT 130.74 439.12 134.79 439.28 ;
      RECT 130.74 439 130.96 439.28 ;
      RECT 130.74 441.04 130.96 441.32 ;
      RECT 130.74 441.04 134.79 441.2 ;
      RECT 130.74 442.52 134.79 442.68 ;
      RECT 130.74 442.4 130.96 442.68 ;
      RECT 130.74 444.44 130.96 444.72 ;
      RECT 130.74 444.44 134.79 444.6 ;
      RECT 130.74 445.92 134.79 446.08 ;
      RECT 130.74 445.8 130.96 446.08 ;
      RECT 130.74 447.84 130.96 448.12 ;
      RECT 130.74 447.84 134.79 448 ;
      RECT 130.74 449.32 134.79 449.48 ;
      RECT 130.74 449.2 130.96 449.48 ;
      RECT 130.74 451.24 130.96 451.52 ;
      RECT 130.74 451.24 134.79 451.4 ;
      RECT 130.74 452.72 134.79 452.88 ;
      RECT 130.74 452.6 130.96 452.88 ;
      RECT 130.74 454.64 130.96 454.92 ;
      RECT 130.74 454.64 134.79 454.8 ;
      RECT 130.74 456.12 134.79 456.28 ;
      RECT 130.74 456 130.96 456.28 ;
      RECT 130.74 458.04 130.96 458.32 ;
      RECT 130.74 458.04 134.79 458.2 ;
      RECT 130.74 459.52 134.79 459.68 ;
      RECT 130.74 459.4 130.96 459.68 ;
      RECT 130.74 461.44 130.96 461.72 ;
      RECT 130.74 461.44 134.79 461.6 ;
      RECT 130.74 462.92 134.79 463.08 ;
      RECT 130.74 462.8 130.96 463.08 ;
      RECT 130.74 464.84 130.96 465.12 ;
      RECT 130.74 464.84 134.79 465 ;
      RECT 130.74 466.32 134.79 466.48 ;
      RECT 130.74 466.2 130.96 466.48 ;
      RECT 130.74 468.24 130.96 468.52 ;
      RECT 130.74 468.24 134.79 468.4 ;
      RECT 130.74 469.72 134.79 469.88 ;
      RECT 130.74 469.6 130.96 469.88 ;
      RECT 130.74 471.64 130.96 471.92 ;
      RECT 130.74 471.64 134.79 471.8 ;
      RECT 130.74 473.12 134.79 473.28 ;
      RECT 130.74 473 130.96 473.28 ;
      RECT 130.74 475.04 130.96 475.32 ;
      RECT 130.74 475.04 134.79 475.2 ;
      RECT 130.74 476.52 134.79 476.68 ;
      RECT 130.74 476.4 130.96 476.68 ;
      RECT 130.74 478.44 130.96 478.72 ;
      RECT 130.74 478.44 134.79 478.6 ;
      RECT 130.74 479.92 134.79 480.08 ;
      RECT 130.74 479.8 130.96 480.08 ;
      RECT 130.74 481.84 130.96 482.12 ;
      RECT 130.74 481.84 134.79 482 ;
      RECT 130.74 483.32 134.79 483.48 ;
      RECT 130.74 483.2 130.96 483.48 ;
      RECT 130.74 485.24 130.96 485.52 ;
      RECT 130.74 485.24 134.79 485.4 ;
      RECT 130.74 486.72 134.79 486.88 ;
      RECT 130.74 486.6 130.96 486.88 ;
      RECT 130.74 488.64 130.96 488.92 ;
      RECT 130.74 488.64 134.79 488.8 ;
      RECT 130.74 490.12 134.79 490.28 ;
      RECT 130.74 490 130.96 490.28 ;
      RECT 130.74 492.04 130.96 492.32 ;
      RECT 130.74 492.04 134.79 492.2 ;
      RECT 130.74 493.52 134.79 493.68 ;
      RECT 130.74 493.4 130.96 493.68 ;
      RECT 130.74 495.44 130.96 495.72 ;
      RECT 130.74 495.44 134.79 495.6 ;
      RECT 130.74 496.92 134.79 497.08 ;
      RECT 130.74 496.8 130.96 497.08 ;
      RECT 130.74 498.84 130.96 499.12 ;
      RECT 130.74 498.84 134.79 499 ;
      RECT 130.74 500.32 134.79 500.48 ;
      RECT 130.74 500.2 130.96 500.48 ;
      RECT 130.74 502.24 130.96 502.52 ;
      RECT 130.74 502.24 134.79 502.4 ;
      RECT 130.74 503.72 134.79 503.88 ;
      RECT 130.74 503.6 130.96 503.88 ;
      RECT 134.15 32.85 134.31 35.75 ;
      RECT 134.31 31.09 134.47 33.01 ;
      RECT 134.31 49.44 134.47 51.3 ;
      RECT 134.15 46.54 134.31 49.6 ;
      RECT 133.73 12.8 134.39 13.06 ;
      RECT 133.73 12.19 133.97 13.06 ;
      RECT 134.15 14.52 134.31 16.86 ;
      RECT 134.02 13.22 134.18 14.84 ;
      RECT 133.75 41.08 133.91 45.17 ;
      RECT 133.75 41.08 134.07 41.24 ;
      RECT 132.93 17.6 133.09 23.81 ;
      RECT 132.45 22.38 133.57 22.54 ;
      RECT 132.93 58.24 133.09 64 ;
      RECT 132.45 59.51 133.57 59.67 ;
      RECT 133.35 27.37 133.51 31.49 ;
      RECT 132.51 27.37 132.67 31.49 ;
      RECT 132.51 27.37 133.51 27.53 ;
      RECT 132.93 24.64 133.09 27.53 ;
      RECT 132.93 54.16 133.09 57.42 ;
      RECT 132.51 54.16 133.51 54.88 ;
      RECT 133.35 50.8 133.51 54.88 ;
      RECT 132.51 50.8 132.67 54.88 ;
      RECT 130.77 55.09 132.03 55.25 ;
      RECT 131.87 49.77 132.03 55.25 ;
      RECT 131.87 49.77 132.75 49.93 ;
      RECT 132.59 32.48 132.75 49.93 ;
      RECT 131.93 45.9 132.75 46.06 ;
      RECT 131.93 36.23 132.75 36.39 ;
      RECT 131.87 32.48 132.75 32.64 ;
      RECT 131.87 27.04 132.03 32.64 ;
      RECT 130.77 27.04 132.03 27.2 ;
      RECT 130.67 26.46 132.69 26.62 ;
      RECT 132.53 25.35 132.69 26.62 ;
      RECT 132.45 22.91 132.61 25.51 ;
      RECT 132.45 56.46 132.61 59.14 ;
      RECT 132.53 55.49 132.69 56.62 ;
      RECT 130.67 55.49 132.69 55.65 ;
      RECT 132.13 25.79 132.37 26.07 ;
      RECT 132.13 21.94 132.29 26.07 ;
      RECT 132.13 21.94 132.41 22.18 ;
      RECT 132.19 15.28 132.35 22.18 ;
      RECT 131.23 15.28 131.39 20.88 ;
      RECT 130.27 15.28 130.43 20.88 ;
      RECT 130.27 17.14 132.35 17.3 ;
      RECT 132.19 59.87 132.35 66.77 ;
      RECT 131.23 61.17 131.39 66.77 ;
      RECT 130.27 61.17 130.43 66.77 ;
      RECT 130.27 64.75 132.35 64.91 ;
      RECT 132.13 59.87 132.41 60.11 ;
      RECT 132.13 56.02 132.29 60.11 ;
      RECT 132.13 56.02 132.37 56.3 ;
      RECT 130.27 35.91 132.35 36.07 ;
      RECT 132.19 32.85 132.35 36.07 ;
      RECT 131.23 27.43 131.39 36.07 ;
      RECT 130.27 32.85 130.43 36.07 ;
      RECT 130.33 27.43 131.39 27.59 ;
      RECT 130.33 23.41 130.49 27.59 ;
      RECT 130.33 26.14 131.49 26.3 ;
      RECT 131.33 25.01 131.49 26.3 ;
      RECT 130.33 25 130.53 26.3 ;
      RECT 131.33 21.38 131.49 23.81 ;
      RECT 130.37 21.38 130.53 23.55 ;
      RECT 130.37 21.38 131.49 21.54 ;
      RECT 130.37 60.51 131.49 60.67 ;
      RECT 131.33 58.24 131.49 60.67 ;
      RECT 130.37 58.5 130.53 60.67 ;
      RECT 130.33 55.81 130.49 58.64 ;
      RECT 131.33 55.81 131.49 57.09 ;
      RECT 130.31 55.81 130.53 57.09 ;
      RECT 130.31 55.81 131.49 55.97 ;
      RECT 130.31 54.64 130.47 57.09 ;
      RECT 130.31 54.64 131.39 54.8 ;
      RECT 131.23 46.22 131.39 54.8 ;
      RECT 132.19 46.22 132.35 49.44 ;
      RECT 130.27 46.22 130.43 49.44 ;
      RECT 130.27 46.22 132.35 46.38 ;
      RECT 131.63 12.8 132.29 13.06 ;
      RECT 132.05 12.19 132.29 13.06 ;
      RECT 132.11 41.08 132.27 45.17 ;
      RECT 131.95 41.08 132.27 41.24 ;
      RECT 121.97 507.88 132.09 508.12 ;
      RECT 114.62 507.74 122.24 507.94 ;
      RECT 121.97 507.38 122.24 508.12 ;
      RECT 114.62 506.28 114.78 507.94 ;
      RECT 114.62 506.28 121.44 506.44 ;
      RECT 120.18 504.68 120.34 506.44 ;
      RECT 118.49 504.68 122.66 504.84 ;
      RECT 119.4 503.72 119.56 504.84 ;
      RECT 119.4 503.72 120.4 503.91 ;
      RECT 131.81 21.06 131.97 26.28 ;
      RECT 130.85 24.37 131.01 25.98 ;
      RECT 130.65 24.37 131.97 24.53 ;
      RECT 130.65 23.67 130.81 24.53 ;
      RECT 130.65 23.67 131.01 23.83 ;
      RECT 130.85 21.7 131.01 23.83 ;
      RECT 130.15 21.06 132.03 21.22 ;
      RECT 130.15 60.83 132.03 60.99 ;
      RECT 131.81 55.81 131.97 60.99 ;
      RECT 130.85 58.22 131.01 60.35 ;
      RECT 130.65 58.22 131.01 58.38 ;
      RECT 130.65 57.25 130.81 58.38 ;
      RECT 130.65 57.25 131.97 57.41 ;
      RECT 130.85 56.13 131.01 57.41 ;
      RECT 131.71 14.52 131.87 16.86 ;
      RECT 131.84 13.22 132 14.84 ;
      RECT 131.71 32.85 131.87 35.75 ;
      RECT 131.55 31.09 131.71 33.01 ;
      RECT 131.55 49.44 131.71 51.3 ;
      RECT 131.71 46.54 131.87 49.6 ;
      RECT 131.63 38.57 131.79 45.17 ;
      RECT 131.33 38.57 131.79 38.73 ;
      RECT 131.33 36.23 131.49 38.73 ;
      RECT 130.97 36.23 131.65 36.39 ;
      RECT 130.85 45.9 131.65 46.06 ;
      RECT 130.85 44.89 131.01 46.06 ;
      RECT 130.83 38.57 130.99 45.17 ;
      RECT 131.23 10.09 131.39 14.2 ;
      RECT 130.33 12.9 131.39 13.06 ;
      RECT 130.33 12.19 130.49 13.06 ;
      RECT 125.55 506.94 130.96 507.15 ;
      RECT 130.76 505.48 130.96 507.15 ;
      RECT 127.34 505.38 127.5 507.15 ;
      RECT 130.75 14.52 130.91 16.86 ;
      RECT 130.62 13.22 130.78 14.84 ;
      RECT 130.75 31.09 130.91 35.75 ;
      RECT 130.65 32.25 130.91 32.53 ;
      RECT 130.71 49.75 130.91 51.3 ;
      RECT 130.75 46.54 130.91 51.3 ;
      RECT 130.31 49.6 130.47 51.7 ;
      RECT 129.87 49.6 130.47 49.76 ;
      RECT 129.87 32.06 130.03 49.76 ;
      RECT 129.87 45.9 130.69 46.06 ;
      RECT 129.87 36.23 130.69 36.39 ;
      RECT 129.87 32.06 130.47 32.22 ;
      RECT 130.31 30.54 130.47 32.22 ;
      RECT 130.35 41.08 130.51 45.17 ;
      RECT 130.35 41.08 130.67 41.24 ;
      RECT 129.52 70.68 130.58 70.84 ;
      RECT 129.52 70.28 129.8 70.84 ;
      RECT 129.52 70.28 130.58 70.44 ;
      RECT 129.52 72.08 130.58 72.24 ;
      RECT 129.52 71.68 129.8 72.24 ;
      RECT 129.52 71.68 130.58 71.84 ;
      RECT 129.52 74.08 130.58 74.24 ;
      RECT 129.52 73.68 129.8 74.24 ;
      RECT 129.52 73.68 130.58 73.84 ;
      RECT 129.52 75.48 130.58 75.64 ;
      RECT 129.52 75.08 129.8 75.64 ;
      RECT 129.52 75.08 130.58 75.24 ;
      RECT 129.52 77.48 130.58 77.64 ;
      RECT 129.52 77.08 129.8 77.64 ;
      RECT 129.52 77.08 130.58 77.24 ;
      RECT 129.52 78.88 130.58 79.04 ;
      RECT 129.52 78.48 129.8 79.04 ;
      RECT 129.52 78.48 130.58 78.64 ;
      RECT 129.52 80.88 130.58 81.04 ;
      RECT 129.52 80.48 129.8 81.04 ;
      RECT 129.52 80.48 130.58 80.64 ;
      RECT 129.52 82.28 130.58 82.44 ;
      RECT 129.52 81.88 129.8 82.44 ;
      RECT 129.52 81.88 130.58 82.04 ;
      RECT 129.52 84.28 130.58 84.44 ;
      RECT 129.52 83.88 129.8 84.44 ;
      RECT 129.52 83.88 130.58 84.04 ;
      RECT 129.52 85.68 130.58 85.84 ;
      RECT 129.52 85.28 129.8 85.84 ;
      RECT 129.52 85.28 130.58 85.44 ;
      RECT 129.52 87.68 130.58 87.84 ;
      RECT 129.52 87.28 129.8 87.84 ;
      RECT 129.52 87.28 130.58 87.44 ;
      RECT 129.52 89.08 130.58 89.24 ;
      RECT 129.52 88.68 129.8 89.24 ;
      RECT 129.52 88.68 130.58 88.84 ;
      RECT 129.52 91.08 130.58 91.24 ;
      RECT 129.52 90.68 129.8 91.24 ;
      RECT 129.52 90.68 130.58 90.84 ;
      RECT 129.52 92.48 130.58 92.64 ;
      RECT 129.52 92.08 129.8 92.64 ;
      RECT 129.52 92.08 130.58 92.24 ;
      RECT 129.52 94.48 130.58 94.64 ;
      RECT 129.52 94.08 129.8 94.64 ;
      RECT 129.52 94.08 130.58 94.24 ;
      RECT 129.52 95.88 130.58 96.04 ;
      RECT 129.52 95.48 129.8 96.04 ;
      RECT 129.52 95.48 130.58 95.64 ;
      RECT 129.52 97.88 130.58 98.04 ;
      RECT 129.52 97.48 129.8 98.04 ;
      RECT 129.52 97.48 130.58 97.64 ;
      RECT 129.52 99.28 130.58 99.44 ;
      RECT 129.52 98.88 129.8 99.44 ;
      RECT 129.52 98.88 130.58 99.04 ;
      RECT 129.52 101.28 130.58 101.44 ;
      RECT 129.52 100.88 129.8 101.44 ;
      RECT 129.52 100.88 130.58 101.04 ;
      RECT 129.52 102.68 130.58 102.84 ;
      RECT 129.52 102.28 129.8 102.84 ;
      RECT 129.52 102.28 130.58 102.44 ;
      RECT 129.52 104.68 130.58 104.84 ;
      RECT 129.52 104.28 129.8 104.84 ;
      RECT 129.52 104.28 130.58 104.44 ;
      RECT 129.52 106.08 130.58 106.24 ;
      RECT 129.52 105.68 129.8 106.24 ;
      RECT 129.52 105.68 130.58 105.84 ;
      RECT 129.52 108.08 130.58 108.24 ;
      RECT 129.52 107.68 129.8 108.24 ;
      RECT 129.52 107.68 130.58 107.84 ;
      RECT 129.52 109.48 130.58 109.64 ;
      RECT 129.52 109.08 129.8 109.64 ;
      RECT 129.52 109.08 130.58 109.24 ;
      RECT 129.52 111.48 130.58 111.64 ;
      RECT 129.52 111.08 129.8 111.64 ;
      RECT 129.52 111.08 130.58 111.24 ;
      RECT 129.52 112.88 130.58 113.04 ;
      RECT 129.52 112.48 129.8 113.04 ;
      RECT 129.52 112.48 130.58 112.64 ;
      RECT 129.52 114.88 130.58 115.04 ;
      RECT 129.52 114.48 129.8 115.04 ;
      RECT 129.52 114.48 130.58 114.64 ;
      RECT 129.52 116.28 130.58 116.44 ;
      RECT 129.52 115.88 129.8 116.44 ;
      RECT 129.52 115.88 130.58 116.04 ;
      RECT 129.52 118.28 130.58 118.44 ;
      RECT 129.52 117.88 129.8 118.44 ;
      RECT 129.52 117.88 130.58 118.04 ;
      RECT 129.52 119.68 130.58 119.84 ;
      RECT 129.52 119.28 129.8 119.84 ;
      RECT 129.52 119.28 130.58 119.44 ;
      RECT 129.52 121.68 130.58 121.84 ;
      RECT 129.52 121.28 129.8 121.84 ;
      RECT 129.52 121.28 130.58 121.44 ;
      RECT 129.52 123.08 130.58 123.24 ;
      RECT 129.52 122.68 129.8 123.24 ;
      RECT 129.52 122.68 130.58 122.84 ;
      RECT 129.52 125.08 130.58 125.24 ;
      RECT 129.52 124.68 129.8 125.24 ;
      RECT 129.52 124.68 130.58 124.84 ;
      RECT 129.52 126.48 130.58 126.64 ;
      RECT 129.52 126.08 129.8 126.64 ;
      RECT 129.52 126.08 130.58 126.24 ;
      RECT 129.52 128.48 130.58 128.64 ;
      RECT 129.52 128.08 129.8 128.64 ;
      RECT 129.52 128.08 130.58 128.24 ;
      RECT 129.52 129.88 130.58 130.04 ;
      RECT 129.52 129.48 129.8 130.04 ;
      RECT 129.52 129.48 130.58 129.64 ;
      RECT 129.52 131.88 130.58 132.04 ;
      RECT 129.52 131.48 129.8 132.04 ;
      RECT 129.52 131.48 130.58 131.64 ;
      RECT 129.52 133.28 130.58 133.44 ;
      RECT 129.52 132.88 129.8 133.44 ;
      RECT 129.52 132.88 130.58 133.04 ;
      RECT 129.52 135.28 130.58 135.44 ;
      RECT 129.52 134.88 129.8 135.44 ;
      RECT 129.52 134.88 130.58 135.04 ;
      RECT 129.52 136.68 130.58 136.84 ;
      RECT 129.52 136.28 129.8 136.84 ;
      RECT 129.52 136.28 130.58 136.44 ;
      RECT 129.52 138.68 130.58 138.84 ;
      RECT 129.52 138.28 129.8 138.84 ;
      RECT 129.52 138.28 130.58 138.44 ;
      RECT 129.52 140.08 130.58 140.24 ;
      RECT 129.52 139.68 129.8 140.24 ;
      RECT 129.52 139.68 130.58 139.84 ;
      RECT 129.52 142.08 130.58 142.24 ;
      RECT 129.52 141.68 129.8 142.24 ;
      RECT 129.52 141.68 130.58 141.84 ;
      RECT 129.52 143.48 130.58 143.64 ;
      RECT 129.52 143.08 129.8 143.64 ;
      RECT 129.52 143.08 130.58 143.24 ;
      RECT 129.52 145.48 130.58 145.64 ;
      RECT 129.52 145.08 129.8 145.64 ;
      RECT 129.52 145.08 130.58 145.24 ;
      RECT 129.52 146.88 130.58 147.04 ;
      RECT 129.52 146.48 129.8 147.04 ;
      RECT 129.52 146.48 130.58 146.64 ;
      RECT 129.52 148.88 130.58 149.04 ;
      RECT 129.52 148.48 129.8 149.04 ;
      RECT 129.52 148.48 130.58 148.64 ;
      RECT 129.52 150.28 130.58 150.44 ;
      RECT 129.52 149.88 129.8 150.44 ;
      RECT 129.52 149.88 130.58 150.04 ;
      RECT 129.52 152.28 130.58 152.44 ;
      RECT 129.52 151.88 129.8 152.44 ;
      RECT 129.52 151.88 130.58 152.04 ;
      RECT 129.52 153.68 130.58 153.84 ;
      RECT 129.52 153.28 129.8 153.84 ;
      RECT 129.52 153.28 130.58 153.44 ;
      RECT 129.52 155.68 130.58 155.84 ;
      RECT 129.52 155.28 129.8 155.84 ;
      RECT 129.52 155.28 130.58 155.44 ;
      RECT 129.52 157.08 130.58 157.24 ;
      RECT 129.52 156.68 129.8 157.24 ;
      RECT 129.52 156.68 130.58 156.84 ;
      RECT 129.52 159.08 130.58 159.24 ;
      RECT 129.52 158.68 129.8 159.24 ;
      RECT 129.52 158.68 130.58 158.84 ;
      RECT 129.52 160.48 130.58 160.64 ;
      RECT 129.52 160.08 129.8 160.64 ;
      RECT 129.52 160.08 130.58 160.24 ;
      RECT 129.52 162.48 130.58 162.64 ;
      RECT 129.52 162.08 129.8 162.64 ;
      RECT 129.52 162.08 130.58 162.24 ;
      RECT 129.52 163.88 130.58 164.04 ;
      RECT 129.52 163.48 129.8 164.04 ;
      RECT 129.52 163.48 130.58 163.64 ;
      RECT 129.52 165.88 130.58 166.04 ;
      RECT 129.52 165.48 129.8 166.04 ;
      RECT 129.52 165.48 130.58 165.64 ;
      RECT 129.52 167.28 130.58 167.44 ;
      RECT 129.52 166.88 129.8 167.44 ;
      RECT 129.52 166.88 130.58 167.04 ;
      RECT 129.52 169.28 130.58 169.44 ;
      RECT 129.52 168.88 129.8 169.44 ;
      RECT 129.52 168.88 130.58 169.04 ;
      RECT 129.52 170.68 130.58 170.84 ;
      RECT 129.52 170.28 129.8 170.84 ;
      RECT 129.52 170.28 130.58 170.44 ;
      RECT 129.52 172.68 130.58 172.84 ;
      RECT 129.52 172.28 129.8 172.84 ;
      RECT 129.52 172.28 130.58 172.44 ;
      RECT 129.52 174.08 130.58 174.24 ;
      RECT 129.52 173.68 129.8 174.24 ;
      RECT 129.52 173.68 130.58 173.84 ;
      RECT 129.52 176.08 130.58 176.24 ;
      RECT 129.52 175.68 129.8 176.24 ;
      RECT 129.52 175.68 130.58 175.84 ;
      RECT 129.52 177.48 130.58 177.64 ;
      RECT 129.52 177.08 129.8 177.64 ;
      RECT 129.52 177.08 130.58 177.24 ;
      RECT 129.52 179.48 130.58 179.64 ;
      RECT 129.52 179.08 129.8 179.64 ;
      RECT 129.52 179.08 130.58 179.24 ;
      RECT 129.52 180.88 130.58 181.04 ;
      RECT 129.52 180.48 129.8 181.04 ;
      RECT 129.52 180.48 130.58 180.64 ;
      RECT 129.52 182.88 130.58 183.04 ;
      RECT 129.52 182.48 129.8 183.04 ;
      RECT 129.52 182.48 130.58 182.64 ;
      RECT 129.52 184.28 130.58 184.44 ;
      RECT 129.52 183.88 129.8 184.44 ;
      RECT 129.52 183.88 130.58 184.04 ;
      RECT 129.52 186.28 130.58 186.44 ;
      RECT 129.52 185.88 129.8 186.44 ;
      RECT 129.52 185.88 130.58 186.04 ;
      RECT 129.52 187.68 130.58 187.84 ;
      RECT 129.52 187.28 129.8 187.84 ;
      RECT 129.52 187.28 130.58 187.44 ;
      RECT 129.52 189.68 130.58 189.84 ;
      RECT 129.52 189.28 129.8 189.84 ;
      RECT 129.52 189.28 130.58 189.44 ;
      RECT 129.52 191.08 130.58 191.24 ;
      RECT 129.52 190.68 129.8 191.24 ;
      RECT 129.52 190.68 130.58 190.84 ;
      RECT 129.52 193.08 130.58 193.24 ;
      RECT 129.52 192.68 129.8 193.24 ;
      RECT 129.52 192.68 130.58 192.84 ;
      RECT 129.52 194.48 130.58 194.64 ;
      RECT 129.52 194.08 129.8 194.64 ;
      RECT 129.52 194.08 130.58 194.24 ;
      RECT 129.52 196.48 130.58 196.64 ;
      RECT 129.52 196.08 129.8 196.64 ;
      RECT 129.52 196.08 130.58 196.24 ;
      RECT 129.52 197.88 130.58 198.04 ;
      RECT 129.52 197.48 129.8 198.04 ;
      RECT 129.52 197.48 130.58 197.64 ;
      RECT 129.52 199.88 130.58 200.04 ;
      RECT 129.52 199.48 129.8 200.04 ;
      RECT 129.52 199.48 130.58 199.64 ;
      RECT 129.52 201.28 130.58 201.44 ;
      RECT 129.52 200.88 129.8 201.44 ;
      RECT 129.52 200.88 130.58 201.04 ;
      RECT 129.52 203.28 130.58 203.44 ;
      RECT 129.52 202.88 129.8 203.44 ;
      RECT 129.52 202.88 130.58 203.04 ;
      RECT 129.52 204.68 130.58 204.84 ;
      RECT 129.52 204.28 129.8 204.84 ;
      RECT 129.52 204.28 130.58 204.44 ;
      RECT 129.52 206.68 130.58 206.84 ;
      RECT 129.52 206.28 129.8 206.84 ;
      RECT 129.52 206.28 130.58 206.44 ;
      RECT 129.52 208.08 130.58 208.24 ;
      RECT 129.52 207.68 129.8 208.24 ;
      RECT 129.52 207.68 130.58 207.84 ;
      RECT 129.52 210.08 130.58 210.24 ;
      RECT 129.52 209.68 129.8 210.24 ;
      RECT 129.52 209.68 130.58 209.84 ;
      RECT 129.52 211.48 130.58 211.64 ;
      RECT 129.52 211.08 129.8 211.64 ;
      RECT 129.52 211.08 130.58 211.24 ;
      RECT 129.52 213.48 130.58 213.64 ;
      RECT 129.52 213.08 129.8 213.64 ;
      RECT 129.52 213.08 130.58 213.24 ;
      RECT 129.52 214.88 130.58 215.04 ;
      RECT 129.52 214.48 129.8 215.04 ;
      RECT 129.52 214.48 130.58 214.64 ;
      RECT 129.52 216.88 130.58 217.04 ;
      RECT 129.52 216.48 129.8 217.04 ;
      RECT 129.52 216.48 130.58 216.64 ;
      RECT 129.52 218.28 130.58 218.44 ;
      RECT 129.52 217.88 129.8 218.44 ;
      RECT 129.52 217.88 130.58 218.04 ;
      RECT 129.52 220.28 130.58 220.44 ;
      RECT 129.52 219.88 129.8 220.44 ;
      RECT 129.52 219.88 130.58 220.04 ;
      RECT 129.52 221.68 130.58 221.84 ;
      RECT 129.52 221.28 129.8 221.84 ;
      RECT 129.52 221.28 130.58 221.44 ;
      RECT 129.52 223.68 130.58 223.84 ;
      RECT 129.52 223.28 129.8 223.84 ;
      RECT 129.52 223.28 130.58 223.44 ;
      RECT 129.52 225.08 130.58 225.24 ;
      RECT 129.52 224.68 129.8 225.24 ;
      RECT 129.52 224.68 130.58 224.84 ;
      RECT 129.52 227.08 130.58 227.24 ;
      RECT 129.52 226.68 129.8 227.24 ;
      RECT 129.52 226.68 130.58 226.84 ;
      RECT 129.52 228.48 130.58 228.64 ;
      RECT 129.52 228.08 129.8 228.64 ;
      RECT 129.52 228.08 130.58 228.24 ;
      RECT 129.52 230.48 130.58 230.64 ;
      RECT 129.52 230.08 129.8 230.64 ;
      RECT 129.52 230.08 130.58 230.24 ;
      RECT 129.52 231.88 130.58 232.04 ;
      RECT 129.52 231.48 129.8 232.04 ;
      RECT 129.52 231.48 130.58 231.64 ;
      RECT 129.52 233.88 130.58 234.04 ;
      RECT 129.52 233.48 129.8 234.04 ;
      RECT 129.52 233.48 130.58 233.64 ;
      RECT 129.52 235.28 130.58 235.44 ;
      RECT 129.52 234.88 129.8 235.44 ;
      RECT 129.52 234.88 130.58 235.04 ;
      RECT 129.52 237.28 130.58 237.44 ;
      RECT 129.52 236.88 129.8 237.44 ;
      RECT 129.52 236.88 130.58 237.04 ;
      RECT 129.52 238.68 130.58 238.84 ;
      RECT 129.52 238.28 129.8 238.84 ;
      RECT 129.52 238.28 130.58 238.44 ;
      RECT 129.52 240.68 130.58 240.84 ;
      RECT 129.52 240.28 129.8 240.84 ;
      RECT 129.52 240.28 130.58 240.44 ;
      RECT 129.52 242.08 130.58 242.24 ;
      RECT 129.52 241.68 129.8 242.24 ;
      RECT 129.52 241.68 130.58 241.84 ;
      RECT 129.52 244.08 130.58 244.24 ;
      RECT 129.52 243.68 129.8 244.24 ;
      RECT 129.52 243.68 130.58 243.84 ;
      RECT 129.52 245.48 130.58 245.64 ;
      RECT 129.52 245.08 129.8 245.64 ;
      RECT 129.52 245.08 130.58 245.24 ;
      RECT 129.52 247.48 130.58 247.64 ;
      RECT 129.52 247.08 129.8 247.64 ;
      RECT 129.52 247.08 130.58 247.24 ;
      RECT 129.52 248.88 130.58 249.04 ;
      RECT 129.52 248.48 129.8 249.04 ;
      RECT 129.52 248.48 130.58 248.64 ;
      RECT 129.52 250.88 130.58 251.04 ;
      RECT 129.52 250.48 129.8 251.04 ;
      RECT 129.52 250.48 130.58 250.64 ;
      RECT 129.52 252.28 130.58 252.44 ;
      RECT 129.52 251.88 129.8 252.44 ;
      RECT 129.52 251.88 130.58 252.04 ;
      RECT 129.52 254.28 130.58 254.44 ;
      RECT 129.52 253.88 129.8 254.44 ;
      RECT 129.52 253.88 130.58 254.04 ;
      RECT 129.52 255.68 130.58 255.84 ;
      RECT 129.52 255.28 129.8 255.84 ;
      RECT 129.52 255.28 130.58 255.44 ;
      RECT 129.52 257.68 130.58 257.84 ;
      RECT 129.52 257.28 129.8 257.84 ;
      RECT 129.52 257.28 130.58 257.44 ;
      RECT 129.52 259.08 130.58 259.24 ;
      RECT 129.52 258.68 129.8 259.24 ;
      RECT 129.52 258.68 130.58 258.84 ;
      RECT 129.52 261.08 130.58 261.24 ;
      RECT 129.52 260.68 129.8 261.24 ;
      RECT 129.52 260.68 130.58 260.84 ;
      RECT 129.52 262.48 130.58 262.64 ;
      RECT 129.52 262.08 129.8 262.64 ;
      RECT 129.52 262.08 130.58 262.24 ;
      RECT 129.52 264.48 130.58 264.64 ;
      RECT 129.52 264.08 129.8 264.64 ;
      RECT 129.52 264.08 130.58 264.24 ;
      RECT 129.52 265.88 130.58 266.04 ;
      RECT 129.52 265.48 129.8 266.04 ;
      RECT 129.52 265.48 130.58 265.64 ;
      RECT 129.52 267.88 130.58 268.04 ;
      RECT 129.52 267.48 129.8 268.04 ;
      RECT 129.52 267.48 130.58 267.64 ;
      RECT 129.52 269.28 130.58 269.44 ;
      RECT 129.52 268.88 129.8 269.44 ;
      RECT 129.52 268.88 130.58 269.04 ;
      RECT 129.52 271.28 130.58 271.44 ;
      RECT 129.52 270.88 129.8 271.44 ;
      RECT 129.52 270.88 130.58 271.04 ;
      RECT 129.52 272.68 130.58 272.84 ;
      RECT 129.52 272.28 129.8 272.84 ;
      RECT 129.52 272.28 130.58 272.44 ;
      RECT 129.52 274.68 130.58 274.84 ;
      RECT 129.52 274.28 129.8 274.84 ;
      RECT 129.52 274.28 130.58 274.44 ;
      RECT 129.52 276.08 130.58 276.24 ;
      RECT 129.52 275.68 129.8 276.24 ;
      RECT 129.52 275.68 130.58 275.84 ;
      RECT 129.52 278.08 130.58 278.24 ;
      RECT 129.52 277.68 129.8 278.24 ;
      RECT 129.52 277.68 130.58 277.84 ;
      RECT 129.52 279.48 130.58 279.64 ;
      RECT 129.52 279.08 129.8 279.64 ;
      RECT 129.52 279.08 130.58 279.24 ;
      RECT 129.52 281.48 130.58 281.64 ;
      RECT 129.52 281.08 129.8 281.64 ;
      RECT 129.52 281.08 130.58 281.24 ;
      RECT 129.52 282.88 130.58 283.04 ;
      RECT 129.52 282.48 129.8 283.04 ;
      RECT 129.52 282.48 130.58 282.64 ;
      RECT 129.52 284.88 130.58 285.04 ;
      RECT 129.52 284.48 129.8 285.04 ;
      RECT 129.52 284.48 130.58 284.64 ;
      RECT 129.52 286.28 130.58 286.44 ;
      RECT 129.52 285.88 129.8 286.44 ;
      RECT 129.52 285.88 130.58 286.04 ;
      RECT 129.52 288.28 130.58 288.44 ;
      RECT 129.52 287.88 129.8 288.44 ;
      RECT 129.52 287.88 130.58 288.04 ;
      RECT 129.52 289.68 130.58 289.84 ;
      RECT 129.52 289.28 129.8 289.84 ;
      RECT 129.52 289.28 130.58 289.44 ;
      RECT 129.52 291.68 130.58 291.84 ;
      RECT 129.52 291.28 129.8 291.84 ;
      RECT 129.52 291.28 130.58 291.44 ;
      RECT 129.52 293.08 130.58 293.24 ;
      RECT 129.52 292.68 129.8 293.24 ;
      RECT 129.52 292.68 130.58 292.84 ;
      RECT 129.52 295.08 130.58 295.24 ;
      RECT 129.52 294.68 129.8 295.24 ;
      RECT 129.52 294.68 130.58 294.84 ;
      RECT 129.52 296.48 130.58 296.64 ;
      RECT 129.52 296.08 129.8 296.64 ;
      RECT 129.52 296.08 130.58 296.24 ;
      RECT 129.52 298.48 130.58 298.64 ;
      RECT 129.52 298.08 129.8 298.64 ;
      RECT 129.52 298.08 130.58 298.24 ;
      RECT 129.52 299.88 130.58 300.04 ;
      RECT 129.52 299.48 129.8 300.04 ;
      RECT 129.52 299.48 130.58 299.64 ;
      RECT 129.52 301.88 130.58 302.04 ;
      RECT 129.52 301.48 129.8 302.04 ;
      RECT 129.52 301.48 130.58 301.64 ;
      RECT 129.52 303.28 130.58 303.44 ;
      RECT 129.52 302.88 129.8 303.44 ;
      RECT 129.52 302.88 130.58 303.04 ;
      RECT 129.52 305.28 130.58 305.44 ;
      RECT 129.52 304.88 129.8 305.44 ;
      RECT 129.52 304.88 130.58 305.04 ;
      RECT 129.52 306.68 130.58 306.84 ;
      RECT 129.52 306.28 129.8 306.84 ;
      RECT 129.52 306.28 130.58 306.44 ;
      RECT 129.52 308.68 130.58 308.84 ;
      RECT 129.52 308.28 129.8 308.84 ;
      RECT 129.52 308.28 130.58 308.44 ;
      RECT 129.52 310.08 130.58 310.24 ;
      RECT 129.52 309.68 129.8 310.24 ;
      RECT 129.52 309.68 130.58 309.84 ;
      RECT 129.52 312.08 130.58 312.24 ;
      RECT 129.52 311.68 129.8 312.24 ;
      RECT 129.52 311.68 130.58 311.84 ;
      RECT 129.52 313.48 130.58 313.64 ;
      RECT 129.52 313.08 129.8 313.64 ;
      RECT 129.52 313.08 130.58 313.24 ;
      RECT 129.52 315.48 130.58 315.64 ;
      RECT 129.52 315.08 129.8 315.64 ;
      RECT 129.52 315.08 130.58 315.24 ;
      RECT 129.52 316.88 130.58 317.04 ;
      RECT 129.52 316.48 129.8 317.04 ;
      RECT 129.52 316.48 130.58 316.64 ;
      RECT 129.52 318.88 130.58 319.04 ;
      RECT 129.52 318.48 129.8 319.04 ;
      RECT 129.52 318.48 130.58 318.64 ;
      RECT 129.52 320.28 130.58 320.44 ;
      RECT 129.52 319.88 129.8 320.44 ;
      RECT 129.52 319.88 130.58 320.04 ;
      RECT 129.52 322.28 130.58 322.44 ;
      RECT 129.52 321.88 129.8 322.44 ;
      RECT 129.52 321.88 130.58 322.04 ;
      RECT 129.52 323.68 130.58 323.84 ;
      RECT 129.52 323.28 129.8 323.84 ;
      RECT 129.52 323.28 130.58 323.44 ;
      RECT 129.52 325.68 130.58 325.84 ;
      RECT 129.52 325.28 129.8 325.84 ;
      RECT 129.52 325.28 130.58 325.44 ;
      RECT 129.52 327.08 130.58 327.24 ;
      RECT 129.52 326.68 129.8 327.24 ;
      RECT 129.52 326.68 130.58 326.84 ;
      RECT 129.52 329.08 130.58 329.24 ;
      RECT 129.52 328.68 129.8 329.24 ;
      RECT 129.52 328.68 130.58 328.84 ;
      RECT 129.52 330.48 130.58 330.64 ;
      RECT 129.52 330.08 129.8 330.64 ;
      RECT 129.52 330.08 130.58 330.24 ;
      RECT 129.52 332.48 130.58 332.64 ;
      RECT 129.52 332.08 129.8 332.64 ;
      RECT 129.52 332.08 130.58 332.24 ;
      RECT 129.52 333.88 130.58 334.04 ;
      RECT 129.52 333.48 129.8 334.04 ;
      RECT 129.52 333.48 130.58 333.64 ;
      RECT 129.52 335.88 130.58 336.04 ;
      RECT 129.52 335.48 129.8 336.04 ;
      RECT 129.52 335.48 130.58 335.64 ;
      RECT 129.52 337.28 130.58 337.44 ;
      RECT 129.52 336.88 129.8 337.44 ;
      RECT 129.52 336.88 130.58 337.04 ;
      RECT 129.52 339.28 130.58 339.44 ;
      RECT 129.52 338.88 129.8 339.44 ;
      RECT 129.52 338.88 130.58 339.04 ;
      RECT 129.52 340.68 130.58 340.84 ;
      RECT 129.52 340.28 129.8 340.84 ;
      RECT 129.52 340.28 130.58 340.44 ;
      RECT 129.52 342.68 130.58 342.84 ;
      RECT 129.52 342.28 129.8 342.84 ;
      RECT 129.52 342.28 130.58 342.44 ;
      RECT 129.52 344.08 130.58 344.24 ;
      RECT 129.52 343.68 129.8 344.24 ;
      RECT 129.52 343.68 130.58 343.84 ;
      RECT 129.52 346.08 130.58 346.24 ;
      RECT 129.52 345.68 129.8 346.24 ;
      RECT 129.52 345.68 130.58 345.84 ;
      RECT 129.52 347.48 130.58 347.64 ;
      RECT 129.52 347.08 129.8 347.64 ;
      RECT 129.52 347.08 130.58 347.24 ;
      RECT 129.52 349.48 130.58 349.64 ;
      RECT 129.52 349.08 129.8 349.64 ;
      RECT 129.52 349.08 130.58 349.24 ;
      RECT 129.52 350.88 130.58 351.04 ;
      RECT 129.52 350.48 129.8 351.04 ;
      RECT 129.52 350.48 130.58 350.64 ;
      RECT 129.52 352.88 130.58 353.04 ;
      RECT 129.52 352.48 129.8 353.04 ;
      RECT 129.52 352.48 130.58 352.64 ;
      RECT 129.52 354.28 130.58 354.44 ;
      RECT 129.52 353.88 129.8 354.44 ;
      RECT 129.52 353.88 130.58 354.04 ;
      RECT 129.52 356.28 130.58 356.44 ;
      RECT 129.52 355.88 129.8 356.44 ;
      RECT 129.52 355.88 130.58 356.04 ;
      RECT 129.52 357.68 130.58 357.84 ;
      RECT 129.52 357.28 129.8 357.84 ;
      RECT 129.52 357.28 130.58 357.44 ;
      RECT 129.52 359.68 130.58 359.84 ;
      RECT 129.52 359.28 129.8 359.84 ;
      RECT 129.52 359.28 130.58 359.44 ;
      RECT 129.52 361.08 130.58 361.24 ;
      RECT 129.52 360.68 129.8 361.24 ;
      RECT 129.52 360.68 130.58 360.84 ;
      RECT 129.52 363.08 130.58 363.24 ;
      RECT 129.52 362.68 129.8 363.24 ;
      RECT 129.52 362.68 130.58 362.84 ;
      RECT 129.52 364.48 130.58 364.64 ;
      RECT 129.52 364.08 129.8 364.64 ;
      RECT 129.52 364.08 130.58 364.24 ;
      RECT 129.52 366.48 130.58 366.64 ;
      RECT 129.52 366.08 129.8 366.64 ;
      RECT 129.52 366.08 130.58 366.24 ;
      RECT 129.52 367.88 130.58 368.04 ;
      RECT 129.52 367.48 129.8 368.04 ;
      RECT 129.52 367.48 130.58 367.64 ;
      RECT 129.52 369.88 130.58 370.04 ;
      RECT 129.52 369.48 129.8 370.04 ;
      RECT 129.52 369.48 130.58 369.64 ;
      RECT 129.52 371.28 130.58 371.44 ;
      RECT 129.52 370.88 129.8 371.44 ;
      RECT 129.52 370.88 130.58 371.04 ;
      RECT 129.52 373.28 130.58 373.44 ;
      RECT 129.52 372.88 129.8 373.44 ;
      RECT 129.52 372.88 130.58 373.04 ;
      RECT 129.52 374.68 130.58 374.84 ;
      RECT 129.52 374.28 129.8 374.84 ;
      RECT 129.52 374.28 130.58 374.44 ;
      RECT 129.52 376.68 130.58 376.84 ;
      RECT 129.52 376.28 129.8 376.84 ;
      RECT 129.52 376.28 130.58 376.44 ;
      RECT 129.52 378.08 130.58 378.24 ;
      RECT 129.52 377.68 129.8 378.24 ;
      RECT 129.52 377.68 130.58 377.84 ;
      RECT 129.52 380.08 130.58 380.24 ;
      RECT 129.52 379.68 129.8 380.24 ;
      RECT 129.52 379.68 130.58 379.84 ;
      RECT 129.52 381.48 130.58 381.64 ;
      RECT 129.52 381.08 129.8 381.64 ;
      RECT 129.52 381.08 130.58 381.24 ;
      RECT 129.52 383.48 130.58 383.64 ;
      RECT 129.52 383.08 129.8 383.64 ;
      RECT 129.52 383.08 130.58 383.24 ;
      RECT 129.52 384.88 130.58 385.04 ;
      RECT 129.52 384.48 129.8 385.04 ;
      RECT 129.52 384.48 130.58 384.64 ;
      RECT 129.52 386.88 130.58 387.04 ;
      RECT 129.52 386.48 129.8 387.04 ;
      RECT 129.52 386.48 130.58 386.64 ;
      RECT 129.52 388.28 130.58 388.44 ;
      RECT 129.52 387.88 129.8 388.44 ;
      RECT 129.52 387.88 130.58 388.04 ;
      RECT 129.52 390.28 130.58 390.44 ;
      RECT 129.52 389.88 129.8 390.44 ;
      RECT 129.52 389.88 130.58 390.04 ;
      RECT 129.52 391.68 130.58 391.84 ;
      RECT 129.52 391.28 129.8 391.84 ;
      RECT 129.52 391.28 130.58 391.44 ;
      RECT 129.52 393.68 130.58 393.84 ;
      RECT 129.52 393.28 129.8 393.84 ;
      RECT 129.52 393.28 130.58 393.44 ;
      RECT 129.52 395.08 130.58 395.24 ;
      RECT 129.52 394.68 129.8 395.24 ;
      RECT 129.52 394.68 130.58 394.84 ;
      RECT 129.52 397.08 130.58 397.24 ;
      RECT 129.52 396.68 129.8 397.24 ;
      RECT 129.52 396.68 130.58 396.84 ;
      RECT 129.52 398.48 130.58 398.64 ;
      RECT 129.52 398.08 129.8 398.64 ;
      RECT 129.52 398.08 130.58 398.24 ;
      RECT 129.52 400.48 130.58 400.64 ;
      RECT 129.52 400.08 129.8 400.64 ;
      RECT 129.52 400.08 130.58 400.24 ;
      RECT 129.52 401.88 130.58 402.04 ;
      RECT 129.52 401.48 129.8 402.04 ;
      RECT 129.52 401.48 130.58 401.64 ;
      RECT 129.52 403.88 130.58 404.04 ;
      RECT 129.52 403.48 129.8 404.04 ;
      RECT 129.52 403.48 130.58 403.64 ;
      RECT 129.52 405.28 130.58 405.44 ;
      RECT 129.52 404.88 129.8 405.44 ;
      RECT 129.52 404.88 130.58 405.04 ;
      RECT 129.52 407.28 130.58 407.44 ;
      RECT 129.52 406.88 129.8 407.44 ;
      RECT 129.52 406.88 130.58 407.04 ;
      RECT 129.52 408.68 130.58 408.84 ;
      RECT 129.52 408.28 129.8 408.84 ;
      RECT 129.52 408.28 130.58 408.44 ;
      RECT 129.52 410.68 130.58 410.84 ;
      RECT 129.52 410.28 129.8 410.84 ;
      RECT 129.52 410.28 130.58 410.44 ;
      RECT 129.52 412.08 130.58 412.24 ;
      RECT 129.52 411.68 129.8 412.24 ;
      RECT 129.52 411.68 130.58 411.84 ;
      RECT 129.52 414.08 130.58 414.24 ;
      RECT 129.52 413.68 129.8 414.24 ;
      RECT 129.52 413.68 130.58 413.84 ;
      RECT 129.52 415.48 130.58 415.64 ;
      RECT 129.52 415.08 129.8 415.64 ;
      RECT 129.52 415.08 130.58 415.24 ;
      RECT 129.52 417.48 130.58 417.64 ;
      RECT 129.52 417.08 129.8 417.64 ;
      RECT 129.52 417.08 130.58 417.24 ;
      RECT 129.52 418.88 130.58 419.04 ;
      RECT 129.52 418.48 129.8 419.04 ;
      RECT 129.52 418.48 130.58 418.64 ;
      RECT 129.52 420.88 130.58 421.04 ;
      RECT 129.52 420.48 129.8 421.04 ;
      RECT 129.52 420.48 130.58 420.64 ;
      RECT 129.52 422.28 130.58 422.44 ;
      RECT 129.52 421.88 129.8 422.44 ;
      RECT 129.52 421.88 130.58 422.04 ;
      RECT 129.52 424.28 130.58 424.44 ;
      RECT 129.52 423.88 129.8 424.44 ;
      RECT 129.52 423.88 130.58 424.04 ;
      RECT 129.52 425.68 130.58 425.84 ;
      RECT 129.52 425.28 129.8 425.84 ;
      RECT 129.52 425.28 130.58 425.44 ;
      RECT 129.52 427.68 130.58 427.84 ;
      RECT 129.52 427.28 129.8 427.84 ;
      RECT 129.52 427.28 130.58 427.44 ;
      RECT 129.52 429.08 130.58 429.24 ;
      RECT 129.52 428.68 129.8 429.24 ;
      RECT 129.52 428.68 130.58 428.84 ;
      RECT 129.52 431.08 130.58 431.24 ;
      RECT 129.52 430.68 129.8 431.24 ;
      RECT 129.52 430.68 130.58 430.84 ;
      RECT 129.52 432.48 130.58 432.64 ;
      RECT 129.52 432.08 129.8 432.64 ;
      RECT 129.52 432.08 130.58 432.24 ;
      RECT 129.52 434.48 130.58 434.64 ;
      RECT 129.52 434.08 129.8 434.64 ;
      RECT 129.52 434.08 130.58 434.24 ;
      RECT 129.52 435.88 130.58 436.04 ;
      RECT 129.52 435.48 129.8 436.04 ;
      RECT 129.52 435.48 130.58 435.64 ;
      RECT 129.52 437.88 130.58 438.04 ;
      RECT 129.52 437.48 129.8 438.04 ;
      RECT 129.52 437.48 130.58 437.64 ;
      RECT 129.52 439.28 130.58 439.44 ;
      RECT 129.52 438.88 129.8 439.44 ;
      RECT 129.52 438.88 130.58 439.04 ;
      RECT 129.52 441.28 130.58 441.44 ;
      RECT 129.52 440.88 129.8 441.44 ;
      RECT 129.52 440.88 130.58 441.04 ;
      RECT 129.52 442.68 130.58 442.84 ;
      RECT 129.52 442.28 129.8 442.84 ;
      RECT 129.52 442.28 130.58 442.44 ;
      RECT 129.52 444.68 130.58 444.84 ;
      RECT 129.52 444.28 129.8 444.84 ;
      RECT 129.52 444.28 130.58 444.44 ;
      RECT 129.52 446.08 130.58 446.24 ;
      RECT 129.52 445.68 129.8 446.24 ;
      RECT 129.52 445.68 130.58 445.84 ;
      RECT 129.52 448.08 130.58 448.24 ;
      RECT 129.52 447.68 129.8 448.24 ;
      RECT 129.52 447.68 130.58 447.84 ;
      RECT 129.52 449.48 130.58 449.64 ;
      RECT 129.52 449.08 129.8 449.64 ;
      RECT 129.52 449.08 130.58 449.24 ;
      RECT 129.52 451.48 130.58 451.64 ;
      RECT 129.52 451.08 129.8 451.64 ;
      RECT 129.52 451.08 130.58 451.24 ;
      RECT 129.52 452.88 130.58 453.04 ;
      RECT 129.52 452.48 129.8 453.04 ;
      RECT 129.52 452.48 130.58 452.64 ;
      RECT 129.52 454.88 130.58 455.04 ;
      RECT 129.52 454.48 129.8 455.04 ;
      RECT 129.52 454.48 130.58 454.64 ;
      RECT 129.52 456.28 130.58 456.44 ;
      RECT 129.52 455.88 129.8 456.44 ;
      RECT 129.52 455.88 130.58 456.04 ;
      RECT 129.52 458.28 130.58 458.44 ;
      RECT 129.52 457.88 129.8 458.44 ;
      RECT 129.52 457.88 130.58 458.04 ;
      RECT 129.52 459.68 130.58 459.84 ;
      RECT 129.52 459.28 129.8 459.84 ;
      RECT 129.52 459.28 130.58 459.44 ;
      RECT 129.52 461.68 130.58 461.84 ;
      RECT 129.52 461.28 129.8 461.84 ;
      RECT 129.52 461.28 130.58 461.44 ;
      RECT 129.52 463.08 130.58 463.24 ;
      RECT 129.52 462.68 129.8 463.24 ;
      RECT 129.52 462.68 130.58 462.84 ;
      RECT 129.52 465.08 130.58 465.24 ;
      RECT 129.52 464.68 129.8 465.24 ;
      RECT 129.52 464.68 130.58 464.84 ;
      RECT 129.52 466.48 130.58 466.64 ;
      RECT 129.52 466.08 129.8 466.64 ;
      RECT 129.52 466.08 130.58 466.24 ;
      RECT 129.52 468.48 130.58 468.64 ;
      RECT 129.52 468.08 129.8 468.64 ;
      RECT 129.52 468.08 130.58 468.24 ;
      RECT 129.52 469.88 130.58 470.04 ;
      RECT 129.52 469.48 129.8 470.04 ;
      RECT 129.52 469.48 130.58 469.64 ;
      RECT 129.52 471.88 130.58 472.04 ;
      RECT 129.52 471.48 129.8 472.04 ;
      RECT 129.52 471.48 130.58 471.64 ;
      RECT 129.52 473.28 130.58 473.44 ;
      RECT 129.52 472.88 129.8 473.44 ;
      RECT 129.52 472.88 130.58 473.04 ;
      RECT 129.52 475.28 130.58 475.44 ;
      RECT 129.52 474.88 129.8 475.44 ;
      RECT 129.52 474.88 130.58 475.04 ;
      RECT 129.52 476.68 130.58 476.84 ;
      RECT 129.52 476.28 129.8 476.84 ;
      RECT 129.52 476.28 130.58 476.44 ;
      RECT 129.52 478.68 130.58 478.84 ;
      RECT 129.52 478.28 129.8 478.84 ;
      RECT 129.52 478.28 130.58 478.44 ;
      RECT 129.52 480.08 130.58 480.24 ;
      RECT 129.52 479.68 129.8 480.24 ;
      RECT 129.52 479.68 130.58 479.84 ;
      RECT 129.52 482.08 130.58 482.24 ;
      RECT 129.52 481.68 129.8 482.24 ;
      RECT 129.52 481.68 130.58 481.84 ;
      RECT 129.52 483.48 130.58 483.64 ;
      RECT 129.52 483.08 129.8 483.64 ;
      RECT 129.52 483.08 130.58 483.24 ;
      RECT 129.52 485.48 130.58 485.64 ;
      RECT 129.52 485.08 129.8 485.64 ;
      RECT 129.52 485.08 130.58 485.24 ;
      RECT 129.52 486.88 130.58 487.04 ;
      RECT 129.52 486.48 129.8 487.04 ;
      RECT 129.52 486.48 130.58 486.64 ;
      RECT 129.52 488.88 130.58 489.04 ;
      RECT 129.52 488.48 129.8 489.04 ;
      RECT 129.52 488.48 130.58 488.64 ;
      RECT 129.52 490.28 130.58 490.44 ;
      RECT 129.52 489.88 129.8 490.44 ;
      RECT 129.52 489.88 130.58 490.04 ;
      RECT 129.52 492.28 130.58 492.44 ;
      RECT 129.52 491.88 129.8 492.44 ;
      RECT 129.52 491.88 130.58 492.04 ;
      RECT 129.52 493.68 130.58 493.84 ;
      RECT 129.52 493.28 129.8 493.84 ;
      RECT 129.52 493.28 130.58 493.44 ;
      RECT 129.52 495.68 130.58 495.84 ;
      RECT 129.52 495.28 129.8 495.84 ;
      RECT 129.52 495.28 130.58 495.44 ;
      RECT 129.52 497.08 130.58 497.24 ;
      RECT 129.52 496.68 129.8 497.24 ;
      RECT 129.52 496.68 130.58 496.84 ;
      RECT 129.52 499.08 130.58 499.24 ;
      RECT 129.52 498.68 129.8 499.24 ;
      RECT 129.52 498.68 130.58 498.84 ;
      RECT 129.52 500.48 130.58 500.64 ;
      RECT 129.52 500.08 129.8 500.64 ;
      RECT 129.52 500.08 130.58 500.24 ;
      RECT 129.52 502.48 130.58 502.64 ;
      RECT 129.52 502.08 129.8 502.64 ;
      RECT 129.52 502.08 130.58 502.24 ;
      RECT 129.52 503.88 130.58 504.04 ;
      RECT 129.52 503.48 129.8 504.04 ;
      RECT 129.52 503.48 130.58 503.64 ;
      RECT 126.63 506.22 127.18 506.5 ;
      RECT 127.02 504.68 127.18 506.5 ;
      RECT 123.49 504.68 130.49 504.84 ;
      RECT 129.53 31.49 129.69 32.02 ;
      RECT 129.07 31.49 130.15 31.65 ;
      RECT 129.99 27.38 130.15 31.65 ;
      RECT 129.07 27.38 129.23 31.65 ;
      RECT 129.07 27.38 130.15 27.54 ;
      RECT 129.53 26.91 129.69 27.54 ;
      RECT 129.07 51.06 130.15 55.29 ;
      RECT 129.53 50.27 129.69 55.29 ;
      RECT 129.74 68.61 130.06 69.01 ;
      RECT 129.27 68.61 130.06 68.77 ;
      RECT 129.89 49.92 130.05 50.9 ;
      RECT 129.17 49.92 129.33 50.9 ;
      RECT 129.17 49.92 130.05 50.08 ;
      RECT 129.53 45.65 129.69 50.08 ;
      RECT 128.75 49.6 128.91 51.7 ;
      RECT 128.75 49.6 129.35 49.76 ;
      RECT 129.19 32.06 129.35 49.76 ;
      RECT 128.53 45.9 129.35 46.06 ;
      RECT 128.53 36.23 129.35 36.39 ;
      RECT 128.75 32.06 129.35 32.22 ;
      RECT 128.75 30.54 128.91 32.22 ;
      RECT 127.25 21.06 127.41 26.28 ;
      RECT 128.21 24.37 128.37 25.98 ;
      RECT 127.25 24.37 128.57 24.53 ;
      RECT 128.41 23.67 128.57 24.53 ;
      RECT 128.21 23.67 128.57 23.83 ;
      RECT 128.21 21.7 128.37 23.83 ;
      RECT 127.19 21.06 129.07 21.22 ;
      RECT 127.19 60.83 129.07 60.99 ;
      RECT 127.25 55.81 127.41 60.99 ;
      RECT 128.21 58.22 128.37 60.35 ;
      RECT 128.21 58.22 128.57 58.38 ;
      RECT 128.41 57.25 128.57 58.38 ;
      RECT 127.25 57.25 128.57 57.41 ;
      RECT 128.21 56.13 128.37 57.41 ;
      RECT 126.85 25.79 127.09 26.07 ;
      RECT 126.93 21.94 127.09 26.07 ;
      RECT 126.81 21.94 127.09 22.18 ;
      RECT 126.87 15.28 127.03 22.18 ;
      RECT 128.79 15.28 128.95 20.88 ;
      RECT 127.83 15.28 127.99 20.88 ;
      RECT 126.87 17.14 128.95 17.3 ;
      RECT 126.87 35.91 128.95 36.07 ;
      RECT 128.79 32.85 128.95 36.07 ;
      RECT 127.83 27.43 127.99 36.07 ;
      RECT 126.87 32.85 127.03 36.07 ;
      RECT 127.83 27.43 128.89 27.59 ;
      RECT 128.73 23.41 128.89 27.59 ;
      RECT 127.73 26.14 128.89 26.3 ;
      RECT 128.69 25 128.89 26.3 ;
      RECT 127.73 25.01 127.89 26.3 ;
      RECT 127.73 21.38 127.89 23.81 ;
      RECT 128.69 21.38 128.85 23.55 ;
      RECT 127.73 21.38 128.85 21.54 ;
      RECT 127.73 60.51 128.85 60.67 ;
      RECT 128.69 58.5 128.85 60.67 ;
      RECT 128.73 55.81 128.85 60.67 ;
      RECT 127.73 58.24 127.89 60.67 ;
      RECT 128.75 54.64 128.89 58.64 ;
      RECT 128.69 55.81 128.91 57.09 ;
      RECT 128.75 54.64 128.91 57.09 ;
      RECT 127.73 55.81 127.89 57.09 ;
      RECT 127.73 55.81 128.91 55.97 ;
      RECT 127.83 54.64 128.91 54.8 ;
      RECT 127.83 46.22 127.99 54.8 ;
      RECT 128.79 46.22 128.95 49.44 ;
      RECT 126.87 46.22 127.03 49.44 ;
      RECT 126.87 46.22 128.95 46.38 ;
      RECT 128.79 61.17 128.95 66.77 ;
      RECT 127.83 61.17 127.99 66.77 ;
      RECT 126.87 59.87 127.03 66.77 ;
      RECT 126.87 64.75 128.95 64.91 ;
      RECT 126.81 59.87 127.09 60.11 ;
      RECT 126.93 56.02 127.09 60.11 ;
      RECT 126.85 56.02 127.09 56.3 ;
      RECT 127.83 10.09 127.99 14.2 ;
      RECT 127.83 12.9 128.89 13.06 ;
      RECT 128.73 12.19 128.89 13.06 ;
      RECT 128.71 41.08 128.87 45.17 ;
      RECT 128.55 41.08 128.87 41.24 ;
      RECT 128.31 14.52 128.47 16.86 ;
      RECT 128.44 13.22 128.6 14.84 ;
      RECT 128.31 31.09 128.47 35.75 ;
      RECT 128.31 32.25 128.57 32.53 ;
      RECT 126.53 26.46 128.55 26.62 ;
      RECT 126.53 25.35 126.69 26.62 ;
      RECT 126.61 22.91 126.77 25.51 ;
      RECT 126.61 56.46 126.77 59.14 ;
      RECT 126.53 55.49 126.69 56.62 ;
      RECT 126.53 55.49 128.55 55.65 ;
      RECT 128.31 49.75 128.51 51.3 ;
      RECT 128.31 46.54 128.47 51.3 ;
      RECT 127.19 55.09 128.45 55.25 ;
      RECT 127.19 49.77 127.35 55.25 ;
      RECT 126.47 49.77 127.35 49.93 ;
      RECT 126.47 32.48 126.63 49.93 ;
      RECT 126.47 45.9 127.29 46.06 ;
      RECT 126.47 36.23 127.29 36.39 ;
      RECT 126.47 32.48 127.35 32.64 ;
      RECT 127.19 27.04 127.35 32.64 ;
      RECT 127.19 27.04 128.45 27.2 ;
      RECT 127.57 45.9 128.37 46.06 ;
      RECT 128.21 44.89 128.37 46.06 ;
      RECT 128.23 38.57 128.39 45.17 ;
      RECT 127.43 38.57 127.59 45.17 ;
      RECT 127.43 38.57 127.89 38.73 ;
      RECT 127.73 36.23 127.89 38.73 ;
      RECT 127.57 36.23 128.25 36.39 ;
      RECT 127.35 32.85 127.51 35.75 ;
      RECT 127.51 31.09 127.67 33.01 ;
      RECT 127.51 49.44 127.67 51.3 ;
      RECT 127.35 46.54 127.51 49.6 ;
      RECT 126.93 12.8 127.59 13.06 ;
      RECT 126.93 12.19 127.17 13.06 ;
      RECT 127.35 14.52 127.51 16.86 ;
      RECT 127.22 13.22 127.38 14.84 ;
      RECT 126.59 70.78 127.34 70.94 ;
      RECT 121.24 70.7 126.75 70.86 ;
      RECT 121.24 70.67 122.02 70.86 ;
      RECT 121.24 71.66 126.75 71.82 ;
      RECT 126.59 71.58 127.34 71.74 ;
      RECT 126.59 74.18 127.34 74.34 ;
      RECT 121.24 74.1 126.75 74.26 ;
      RECT 121.24 75.06 122.02 75.25 ;
      RECT 121.24 75.06 126.75 75.22 ;
      RECT 126.59 74.98 127.34 75.14 ;
      RECT 126.59 77.58 127.34 77.74 ;
      RECT 121.24 77.5 126.75 77.66 ;
      RECT 121.24 77.47 122.02 77.66 ;
      RECT 121.24 78.46 126.75 78.62 ;
      RECT 126.59 78.38 127.34 78.54 ;
      RECT 126.59 80.98 127.34 81.14 ;
      RECT 121.24 80.9 126.75 81.06 ;
      RECT 121.24 81.86 122.02 82.05 ;
      RECT 121.24 81.86 126.75 82.02 ;
      RECT 126.59 81.78 127.34 81.94 ;
      RECT 126.59 84.38 127.34 84.54 ;
      RECT 121.24 84.3 126.75 84.46 ;
      RECT 121.24 84.27 122.02 84.46 ;
      RECT 121.24 85.26 126.75 85.42 ;
      RECT 126.59 85.18 127.34 85.34 ;
      RECT 126.59 87.78 127.34 87.94 ;
      RECT 121.24 87.7 126.75 87.86 ;
      RECT 121.24 88.66 122.02 88.85 ;
      RECT 121.24 88.66 126.75 88.82 ;
      RECT 126.59 88.58 127.34 88.74 ;
      RECT 126.59 91.18 127.34 91.34 ;
      RECT 121.24 91.1 126.75 91.26 ;
      RECT 121.24 91.07 122.02 91.26 ;
      RECT 121.24 92.06 126.75 92.22 ;
      RECT 126.59 91.98 127.34 92.14 ;
      RECT 126.59 94.58 127.34 94.74 ;
      RECT 121.24 94.5 126.75 94.66 ;
      RECT 121.24 95.46 122.02 95.65 ;
      RECT 121.24 95.46 126.75 95.62 ;
      RECT 126.59 95.38 127.34 95.54 ;
      RECT 126.59 97.98 127.34 98.14 ;
      RECT 121.24 97.9 126.75 98.06 ;
      RECT 121.24 97.87 122.02 98.06 ;
      RECT 121.24 98.86 126.75 99.02 ;
      RECT 126.59 98.78 127.34 98.94 ;
      RECT 126.59 101.38 127.34 101.54 ;
      RECT 121.24 101.3 126.75 101.46 ;
      RECT 121.24 102.26 122.02 102.45 ;
      RECT 121.24 102.26 126.75 102.42 ;
      RECT 126.59 102.18 127.34 102.34 ;
      RECT 126.59 104.78 127.34 104.94 ;
      RECT 121.24 104.7 126.75 104.86 ;
      RECT 121.24 104.67 122.02 104.86 ;
      RECT 121.24 105.66 126.75 105.82 ;
      RECT 126.59 105.58 127.34 105.74 ;
      RECT 126.59 108.18 127.34 108.34 ;
      RECT 121.24 108.1 126.75 108.26 ;
      RECT 121.24 109.06 122.02 109.25 ;
      RECT 121.24 109.06 126.75 109.22 ;
      RECT 126.59 108.98 127.34 109.14 ;
      RECT 126.59 111.58 127.34 111.74 ;
      RECT 121.24 111.5 126.75 111.66 ;
      RECT 121.24 111.47 122.02 111.66 ;
      RECT 121.24 112.46 126.75 112.62 ;
      RECT 126.59 112.38 127.34 112.54 ;
      RECT 126.59 114.98 127.34 115.14 ;
      RECT 121.24 114.9 126.75 115.06 ;
      RECT 121.24 115.86 122.02 116.05 ;
      RECT 121.24 115.86 126.75 116.02 ;
      RECT 126.59 115.78 127.34 115.94 ;
      RECT 126.59 118.38 127.34 118.54 ;
      RECT 121.24 118.3 126.75 118.46 ;
      RECT 121.24 118.27 122.02 118.46 ;
      RECT 121.24 119.26 126.75 119.42 ;
      RECT 126.59 119.18 127.34 119.34 ;
      RECT 126.59 121.78 127.34 121.94 ;
      RECT 121.24 121.7 126.75 121.86 ;
      RECT 121.24 122.66 122.02 122.85 ;
      RECT 121.24 122.66 126.75 122.82 ;
      RECT 126.59 122.58 127.34 122.74 ;
      RECT 126.59 125.18 127.34 125.34 ;
      RECT 121.24 125.1 126.75 125.26 ;
      RECT 121.24 125.07 122.02 125.26 ;
      RECT 121.24 126.06 126.75 126.22 ;
      RECT 126.59 125.98 127.34 126.14 ;
      RECT 126.59 128.58 127.34 128.74 ;
      RECT 121.24 128.5 126.75 128.66 ;
      RECT 121.24 129.46 122.02 129.65 ;
      RECT 121.24 129.46 126.75 129.62 ;
      RECT 126.59 129.38 127.34 129.54 ;
      RECT 126.59 131.98 127.34 132.14 ;
      RECT 121.24 131.9 126.75 132.06 ;
      RECT 121.24 131.87 122.02 132.06 ;
      RECT 121.24 132.86 126.75 133.02 ;
      RECT 126.59 132.78 127.34 132.94 ;
      RECT 126.59 135.38 127.34 135.54 ;
      RECT 121.24 135.3 126.75 135.46 ;
      RECT 121.24 136.26 122.02 136.45 ;
      RECT 121.24 136.26 126.75 136.42 ;
      RECT 126.59 136.18 127.34 136.34 ;
      RECT 126.59 138.78 127.34 138.94 ;
      RECT 121.24 138.7 126.75 138.86 ;
      RECT 121.24 138.67 122.02 138.86 ;
      RECT 121.24 139.66 126.75 139.82 ;
      RECT 126.59 139.58 127.34 139.74 ;
      RECT 126.59 142.18 127.34 142.34 ;
      RECT 121.24 142.1 126.75 142.26 ;
      RECT 121.24 143.06 122.02 143.25 ;
      RECT 121.24 143.06 126.75 143.22 ;
      RECT 126.59 142.98 127.34 143.14 ;
      RECT 126.59 145.58 127.34 145.74 ;
      RECT 121.24 145.5 126.75 145.66 ;
      RECT 121.24 145.47 122.02 145.66 ;
      RECT 121.24 146.46 126.75 146.62 ;
      RECT 126.59 146.38 127.34 146.54 ;
      RECT 126.59 148.98 127.34 149.14 ;
      RECT 121.24 148.9 126.75 149.06 ;
      RECT 121.24 149.86 122.02 150.05 ;
      RECT 121.24 149.86 126.75 150.02 ;
      RECT 126.59 149.78 127.34 149.94 ;
      RECT 126.59 152.38 127.34 152.54 ;
      RECT 121.24 152.3 126.75 152.46 ;
      RECT 121.24 152.27 122.02 152.46 ;
      RECT 121.24 153.26 126.75 153.42 ;
      RECT 126.59 153.18 127.34 153.34 ;
      RECT 126.59 155.78 127.34 155.94 ;
      RECT 121.24 155.7 126.75 155.86 ;
      RECT 121.24 156.66 122.02 156.85 ;
      RECT 121.24 156.66 126.75 156.82 ;
      RECT 126.59 156.58 127.34 156.74 ;
      RECT 126.59 159.18 127.34 159.34 ;
      RECT 121.24 159.1 126.75 159.26 ;
      RECT 121.24 159.07 122.02 159.26 ;
      RECT 121.24 160.06 126.75 160.22 ;
      RECT 126.59 159.98 127.34 160.14 ;
      RECT 126.59 162.58 127.34 162.74 ;
      RECT 121.24 162.5 126.75 162.66 ;
      RECT 121.24 163.46 122.02 163.65 ;
      RECT 121.24 163.46 126.75 163.62 ;
      RECT 126.59 163.38 127.34 163.54 ;
      RECT 126.59 165.98 127.34 166.14 ;
      RECT 121.24 165.9 126.75 166.06 ;
      RECT 121.24 165.87 122.02 166.06 ;
      RECT 121.24 166.86 126.75 167.02 ;
      RECT 126.59 166.78 127.34 166.94 ;
      RECT 126.59 169.38 127.34 169.54 ;
      RECT 121.24 169.3 126.75 169.46 ;
      RECT 121.24 170.26 122.02 170.45 ;
      RECT 121.24 170.26 126.75 170.42 ;
      RECT 126.59 170.18 127.34 170.34 ;
      RECT 126.59 172.78 127.34 172.94 ;
      RECT 121.24 172.7 126.75 172.86 ;
      RECT 121.24 172.67 122.02 172.86 ;
      RECT 121.24 173.66 126.75 173.82 ;
      RECT 126.59 173.58 127.34 173.74 ;
      RECT 126.59 176.18 127.34 176.34 ;
      RECT 121.24 176.1 126.75 176.26 ;
      RECT 121.24 177.06 122.02 177.25 ;
      RECT 121.24 177.06 126.75 177.22 ;
      RECT 126.59 176.98 127.34 177.14 ;
      RECT 126.59 179.58 127.34 179.74 ;
      RECT 121.24 179.5 126.75 179.66 ;
      RECT 121.24 179.47 122.02 179.66 ;
      RECT 121.24 180.46 126.75 180.62 ;
      RECT 126.59 180.38 127.34 180.54 ;
      RECT 126.59 182.98 127.34 183.14 ;
      RECT 121.24 182.9 126.75 183.06 ;
      RECT 121.24 183.86 122.02 184.05 ;
      RECT 121.24 183.86 126.75 184.02 ;
      RECT 126.59 183.78 127.34 183.94 ;
      RECT 126.59 186.38 127.34 186.54 ;
      RECT 121.24 186.3 126.75 186.46 ;
      RECT 121.24 186.27 122.02 186.46 ;
      RECT 121.24 187.26 126.75 187.42 ;
      RECT 126.59 187.18 127.34 187.34 ;
      RECT 126.59 189.78 127.34 189.94 ;
      RECT 121.24 189.7 126.75 189.86 ;
      RECT 121.24 190.66 122.02 190.85 ;
      RECT 121.24 190.66 126.75 190.82 ;
      RECT 126.59 190.58 127.34 190.74 ;
      RECT 126.59 193.18 127.34 193.34 ;
      RECT 121.24 193.1 126.75 193.26 ;
      RECT 121.24 193.07 122.02 193.26 ;
      RECT 121.24 194.06 126.75 194.22 ;
      RECT 126.59 193.98 127.34 194.14 ;
      RECT 126.59 196.58 127.34 196.74 ;
      RECT 121.24 196.5 126.75 196.66 ;
      RECT 121.24 197.46 122.02 197.65 ;
      RECT 121.24 197.46 126.75 197.62 ;
      RECT 126.59 197.38 127.34 197.54 ;
      RECT 126.59 199.98 127.34 200.14 ;
      RECT 121.24 199.9 126.75 200.06 ;
      RECT 121.24 199.87 122.02 200.06 ;
      RECT 121.24 200.86 126.75 201.02 ;
      RECT 126.59 200.78 127.34 200.94 ;
      RECT 126.59 203.38 127.34 203.54 ;
      RECT 121.24 203.3 126.75 203.46 ;
      RECT 121.24 204.26 122.02 204.45 ;
      RECT 121.24 204.26 126.75 204.42 ;
      RECT 126.59 204.18 127.34 204.34 ;
      RECT 126.59 206.78 127.34 206.94 ;
      RECT 121.24 206.7 126.75 206.86 ;
      RECT 121.24 206.67 122.02 206.86 ;
      RECT 121.24 207.66 126.75 207.82 ;
      RECT 126.59 207.58 127.34 207.74 ;
      RECT 126.59 210.18 127.34 210.34 ;
      RECT 121.24 210.1 126.75 210.26 ;
      RECT 121.24 211.06 122.02 211.25 ;
      RECT 121.24 211.06 126.75 211.22 ;
      RECT 126.59 210.98 127.34 211.14 ;
      RECT 126.59 213.58 127.34 213.74 ;
      RECT 121.24 213.5 126.75 213.66 ;
      RECT 121.24 213.47 122.02 213.66 ;
      RECT 121.24 214.46 126.75 214.62 ;
      RECT 126.59 214.38 127.34 214.54 ;
      RECT 126.59 216.98 127.34 217.14 ;
      RECT 121.24 216.9 126.75 217.06 ;
      RECT 121.24 217.86 122.02 218.05 ;
      RECT 121.24 217.86 126.75 218.02 ;
      RECT 126.59 217.78 127.34 217.94 ;
      RECT 126.59 220.38 127.34 220.54 ;
      RECT 121.24 220.3 126.75 220.46 ;
      RECT 121.24 220.27 122.02 220.46 ;
      RECT 121.24 221.26 126.75 221.42 ;
      RECT 126.59 221.18 127.34 221.34 ;
      RECT 126.59 223.78 127.34 223.94 ;
      RECT 121.24 223.7 126.75 223.86 ;
      RECT 121.24 224.66 122.02 224.85 ;
      RECT 121.24 224.66 126.75 224.82 ;
      RECT 126.59 224.58 127.34 224.74 ;
      RECT 126.59 227.18 127.34 227.34 ;
      RECT 121.24 227.1 126.75 227.26 ;
      RECT 121.24 227.07 122.02 227.26 ;
      RECT 121.24 228.06 126.75 228.22 ;
      RECT 126.59 227.98 127.34 228.14 ;
      RECT 126.59 230.58 127.34 230.74 ;
      RECT 121.24 230.5 126.75 230.66 ;
      RECT 121.24 231.46 122.02 231.65 ;
      RECT 121.24 231.46 126.75 231.62 ;
      RECT 126.59 231.38 127.34 231.54 ;
      RECT 126.59 233.98 127.34 234.14 ;
      RECT 121.24 233.9 126.75 234.06 ;
      RECT 121.24 233.87 122.02 234.06 ;
      RECT 121.24 234.86 126.75 235.02 ;
      RECT 126.59 234.78 127.34 234.94 ;
      RECT 126.59 237.38 127.34 237.54 ;
      RECT 121.24 237.3 126.75 237.46 ;
      RECT 121.24 238.26 122.02 238.45 ;
      RECT 121.24 238.26 126.75 238.42 ;
      RECT 126.59 238.18 127.34 238.34 ;
      RECT 126.59 240.78 127.34 240.94 ;
      RECT 121.24 240.7 126.75 240.86 ;
      RECT 121.24 240.67 122.02 240.86 ;
      RECT 121.24 241.66 126.75 241.82 ;
      RECT 126.59 241.58 127.34 241.74 ;
      RECT 126.59 244.18 127.34 244.34 ;
      RECT 121.24 244.1 126.75 244.26 ;
      RECT 121.24 245.06 122.02 245.25 ;
      RECT 121.24 245.06 126.75 245.22 ;
      RECT 126.59 244.98 127.34 245.14 ;
      RECT 126.59 247.58 127.34 247.74 ;
      RECT 121.24 247.5 126.75 247.66 ;
      RECT 121.24 247.47 122.02 247.66 ;
      RECT 121.24 248.46 126.75 248.62 ;
      RECT 126.59 248.38 127.34 248.54 ;
      RECT 126.59 250.98 127.34 251.14 ;
      RECT 121.24 250.9 126.75 251.06 ;
      RECT 121.24 251.86 122.02 252.05 ;
      RECT 121.24 251.86 126.75 252.02 ;
      RECT 126.59 251.78 127.34 251.94 ;
      RECT 126.59 254.38 127.34 254.54 ;
      RECT 121.24 254.3 126.75 254.46 ;
      RECT 121.24 254.27 122.02 254.46 ;
      RECT 121.24 255.26 126.75 255.42 ;
      RECT 126.59 255.18 127.34 255.34 ;
      RECT 126.59 257.78 127.34 257.94 ;
      RECT 121.24 257.7 126.75 257.86 ;
      RECT 121.24 258.66 122.02 258.85 ;
      RECT 121.24 258.66 126.75 258.82 ;
      RECT 126.59 258.58 127.34 258.74 ;
      RECT 126.59 261.18 127.34 261.34 ;
      RECT 121.24 261.1 126.75 261.26 ;
      RECT 121.24 261.07 122.02 261.26 ;
      RECT 121.24 262.06 126.75 262.22 ;
      RECT 126.59 261.98 127.34 262.14 ;
      RECT 126.59 264.58 127.34 264.74 ;
      RECT 121.24 264.5 126.75 264.66 ;
      RECT 121.24 265.46 122.02 265.65 ;
      RECT 121.24 265.46 126.75 265.62 ;
      RECT 126.59 265.38 127.34 265.54 ;
      RECT 126.59 267.98 127.34 268.14 ;
      RECT 121.24 267.9 126.75 268.06 ;
      RECT 121.24 267.87 122.02 268.06 ;
      RECT 121.24 268.86 126.75 269.02 ;
      RECT 126.59 268.78 127.34 268.94 ;
      RECT 126.59 271.38 127.34 271.54 ;
      RECT 121.24 271.3 126.75 271.46 ;
      RECT 121.24 272.26 122.02 272.45 ;
      RECT 121.24 272.26 126.75 272.42 ;
      RECT 126.59 272.18 127.34 272.34 ;
      RECT 126.59 274.78 127.34 274.94 ;
      RECT 121.24 274.7 126.75 274.86 ;
      RECT 121.24 274.67 122.02 274.86 ;
      RECT 121.24 275.66 126.75 275.82 ;
      RECT 126.59 275.58 127.34 275.74 ;
      RECT 126.59 278.18 127.34 278.34 ;
      RECT 121.24 278.1 126.75 278.26 ;
      RECT 121.24 279.06 122.02 279.25 ;
      RECT 121.24 279.06 126.75 279.22 ;
      RECT 126.59 278.98 127.34 279.14 ;
      RECT 126.59 281.58 127.34 281.74 ;
      RECT 121.24 281.5 126.75 281.66 ;
      RECT 121.24 281.47 122.02 281.66 ;
      RECT 121.24 282.46 126.75 282.62 ;
      RECT 126.59 282.38 127.34 282.54 ;
      RECT 126.59 284.98 127.34 285.14 ;
      RECT 121.24 284.9 126.75 285.06 ;
      RECT 121.24 285.86 122.02 286.05 ;
      RECT 121.24 285.86 126.75 286.02 ;
      RECT 126.59 285.78 127.34 285.94 ;
      RECT 126.59 288.38 127.34 288.54 ;
      RECT 121.24 288.3 126.75 288.46 ;
      RECT 121.24 288.27 122.02 288.46 ;
      RECT 121.24 289.26 126.75 289.42 ;
      RECT 126.59 289.18 127.34 289.34 ;
      RECT 126.59 291.78 127.34 291.94 ;
      RECT 121.24 291.7 126.75 291.86 ;
      RECT 121.24 292.66 122.02 292.85 ;
      RECT 121.24 292.66 126.75 292.82 ;
      RECT 126.59 292.58 127.34 292.74 ;
      RECT 126.59 295.18 127.34 295.34 ;
      RECT 121.24 295.1 126.75 295.26 ;
      RECT 121.24 295.07 122.02 295.26 ;
      RECT 121.24 296.06 126.75 296.22 ;
      RECT 126.59 295.98 127.34 296.14 ;
      RECT 126.59 298.58 127.34 298.74 ;
      RECT 121.24 298.5 126.75 298.66 ;
      RECT 121.24 299.46 122.02 299.65 ;
      RECT 121.24 299.46 126.75 299.62 ;
      RECT 126.59 299.38 127.34 299.54 ;
      RECT 126.59 301.98 127.34 302.14 ;
      RECT 121.24 301.9 126.75 302.06 ;
      RECT 121.24 301.87 122.02 302.06 ;
      RECT 121.24 302.86 126.75 303.02 ;
      RECT 126.59 302.78 127.34 302.94 ;
      RECT 126.59 305.38 127.34 305.54 ;
      RECT 121.24 305.3 126.75 305.46 ;
      RECT 121.24 306.26 122.02 306.45 ;
      RECT 121.24 306.26 126.75 306.42 ;
      RECT 126.59 306.18 127.34 306.34 ;
      RECT 126.59 308.78 127.34 308.94 ;
      RECT 121.24 308.7 126.75 308.86 ;
      RECT 121.24 308.67 122.02 308.86 ;
      RECT 121.24 309.66 126.75 309.82 ;
      RECT 126.59 309.58 127.34 309.74 ;
      RECT 126.59 312.18 127.34 312.34 ;
      RECT 121.24 312.1 126.75 312.26 ;
      RECT 121.24 313.06 122.02 313.25 ;
      RECT 121.24 313.06 126.75 313.22 ;
      RECT 126.59 312.98 127.34 313.14 ;
      RECT 126.59 315.58 127.34 315.74 ;
      RECT 121.24 315.5 126.75 315.66 ;
      RECT 121.24 315.47 122.02 315.66 ;
      RECT 121.24 316.46 126.75 316.62 ;
      RECT 126.59 316.38 127.34 316.54 ;
      RECT 126.59 318.98 127.34 319.14 ;
      RECT 121.24 318.9 126.75 319.06 ;
      RECT 121.24 319.86 122.02 320.05 ;
      RECT 121.24 319.86 126.75 320.02 ;
      RECT 126.59 319.78 127.34 319.94 ;
      RECT 126.59 322.38 127.34 322.54 ;
      RECT 121.24 322.3 126.75 322.46 ;
      RECT 121.24 322.27 122.02 322.46 ;
      RECT 121.24 323.26 126.75 323.42 ;
      RECT 126.59 323.18 127.34 323.34 ;
      RECT 126.59 325.78 127.34 325.94 ;
      RECT 121.24 325.7 126.75 325.86 ;
      RECT 121.24 326.66 122.02 326.85 ;
      RECT 121.24 326.66 126.75 326.82 ;
      RECT 126.59 326.58 127.34 326.74 ;
      RECT 126.59 329.18 127.34 329.34 ;
      RECT 121.24 329.1 126.75 329.26 ;
      RECT 121.24 329.07 122.02 329.26 ;
      RECT 121.24 330.06 126.75 330.22 ;
      RECT 126.59 329.98 127.34 330.14 ;
      RECT 126.59 332.58 127.34 332.74 ;
      RECT 121.24 332.5 126.75 332.66 ;
      RECT 121.24 333.46 122.02 333.65 ;
      RECT 121.24 333.46 126.75 333.62 ;
      RECT 126.59 333.38 127.34 333.54 ;
      RECT 126.59 335.98 127.34 336.14 ;
      RECT 121.24 335.9 126.75 336.06 ;
      RECT 121.24 335.87 122.02 336.06 ;
      RECT 121.24 336.86 126.75 337.02 ;
      RECT 126.59 336.78 127.34 336.94 ;
      RECT 126.59 339.38 127.34 339.54 ;
      RECT 121.24 339.3 126.75 339.46 ;
      RECT 121.24 340.26 122.02 340.45 ;
      RECT 121.24 340.26 126.75 340.42 ;
      RECT 126.59 340.18 127.34 340.34 ;
      RECT 126.59 342.78 127.34 342.94 ;
      RECT 121.24 342.7 126.75 342.86 ;
      RECT 121.24 342.67 122.02 342.86 ;
      RECT 121.24 343.66 126.75 343.82 ;
      RECT 126.59 343.58 127.34 343.74 ;
      RECT 126.59 346.18 127.34 346.34 ;
      RECT 121.24 346.1 126.75 346.26 ;
      RECT 121.24 347.06 122.02 347.25 ;
      RECT 121.24 347.06 126.75 347.22 ;
      RECT 126.59 346.98 127.34 347.14 ;
      RECT 126.59 349.58 127.34 349.74 ;
      RECT 121.24 349.5 126.75 349.66 ;
      RECT 121.24 349.47 122.02 349.66 ;
      RECT 121.24 350.46 126.75 350.62 ;
      RECT 126.59 350.38 127.34 350.54 ;
      RECT 126.59 352.98 127.34 353.14 ;
      RECT 121.24 352.9 126.75 353.06 ;
      RECT 121.24 353.86 122.02 354.05 ;
      RECT 121.24 353.86 126.75 354.02 ;
      RECT 126.59 353.78 127.34 353.94 ;
      RECT 126.59 356.38 127.34 356.54 ;
      RECT 121.24 356.3 126.75 356.46 ;
      RECT 121.24 356.27 122.02 356.46 ;
      RECT 121.24 357.26 126.75 357.42 ;
      RECT 126.59 357.18 127.34 357.34 ;
      RECT 126.59 359.78 127.34 359.94 ;
      RECT 121.24 359.7 126.75 359.86 ;
      RECT 121.24 360.66 122.02 360.85 ;
      RECT 121.24 360.66 126.75 360.82 ;
      RECT 126.59 360.58 127.34 360.74 ;
      RECT 126.59 363.18 127.34 363.34 ;
      RECT 121.24 363.1 126.75 363.26 ;
      RECT 121.24 363.07 122.02 363.26 ;
      RECT 121.24 364.06 126.75 364.22 ;
      RECT 126.59 363.98 127.34 364.14 ;
      RECT 126.59 366.58 127.34 366.74 ;
      RECT 121.24 366.5 126.75 366.66 ;
      RECT 121.24 367.46 122.02 367.65 ;
      RECT 121.24 367.46 126.75 367.62 ;
      RECT 126.59 367.38 127.34 367.54 ;
      RECT 126.59 369.98 127.34 370.14 ;
      RECT 121.24 369.9 126.75 370.06 ;
      RECT 121.24 369.87 122.02 370.06 ;
      RECT 121.24 370.86 126.75 371.02 ;
      RECT 126.59 370.78 127.34 370.94 ;
      RECT 126.59 373.38 127.34 373.54 ;
      RECT 121.24 373.3 126.75 373.46 ;
      RECT 121.24 374.26 122.02 374.45 ;
      RECT 121.24 374.26 126.75 374.42 ;
      RECT 126.59 374.18 127.34 374.34 ;
      RECT 126.59 376.78 127.34 376.94 ;
      RECT 121.24 376.7 126.75 376.86 ;
      RECT 121.24 376.67 122.02 376.86 ;
      RECT 121.24 377.66 126.75 377.82 ;
      RECT 126.59 377.58 127.34 377.74 ;
      RECT 126.59 380.18 127.34 380.34 ;
      RECT 121.24 380.1 126.75 380.26 ;
      RECT 121.24 381.06 122.02 381.25 ;
      RECT 121.24 381.06 126.75 381.22 ;
      RECT 126.59 380.98 127.34 381.14 ;
      RECT 126.59 383.58 127.34 383.74 ;
      RECT 121.24 383.5 126.75 383.66 ;
      RECT 121.24 383.47 122.02 383.66 ;
      RECT 121.24 384.46 126.75 384.62 ;
      RECT 126.59 384.38 127.34 384.54 ;
      RECT 126.59 386.98 127.34 387.14 ;
      RECT 121.24 386.9 126.75 387.06 ;
      RECT 121.24 387.86 122.02 388.05 ;
      RECT 121.24 387.86 126.75 388.02 ;
      RECT 126.59 387.78 127.34 387.94 ;
      RECT 126.59 390.38 127.34 390.54 ;
      RECT 121.24 390.3 126.75 390.46 ;
      RECT 121.24 390.27 122.02 390.46 ;
      RECT 121.24 391.26 126.75 391.42 ;
      RECT 126.59 391.18 127.34 391.34 ;
      RECT 126.59 393.78 127.34 393.94 ;
      RECT 121.24 393.7 126.75 393.86 ;
      RECT 121.24 394.66 122.02 394.85 ;
      RECT 121.24 394.66 126.75 394.82 ;
      RECT 126.59 394.58 127.34 394.74 ;
      RECT 126.59 397.18 127.34 397.34 ;
      RECT 121.24 397.1 126.75 397.26 ;
      RECT 121.24 397.07 122.02 397.26 ;
      RECT 121.24 398.06 126.75 398.22 ;
      RECT 126.59 397.98 127.34 398.14 ;
      RECT 126.59 400.58 127.34 400.74 ;
      RECT 121.24 400.5 126.75 400.66 ;
      RECT 121.24 401.46 122.02 401.65 ;
      RECT 121.24 401.46 126.75 401.62 ;
      RECT 126.59 401.38 127.34 401.54 ;
      RECT 126.59 403.98 127.34 404.14 ;
      RECT 121.24 403.9 126.75 404.06 ;
      RECT 121.24 403.87 122.02 404.06 ;
      RECT 121.24 404.86 126.75 405.02 ;
      RECT 126.59 404.78 127.34 404.94 ;
      RECT 126.59 407.38 127.34 407.54 ;
      RECT 121.24 407.3 126.75 407.46 ;
      RECT 121.24 408.26 122.02 408.45 ;
      RECT 121.24 408.26 126.75 408.42 ;
      RECT 126.59 408.18 127.34 408.34 ;
      RECT 126.59 410.78 127.34 410.94 ;
      RECT 121.24 410.7 126.75 410.86 ;
      RECT 121.24 410.67 122.02 410.86 ;
      RECT 121.24 411.66 126.75 411.82 ;
      RECT 126.59 411.58 127.34 411.74 ;
      RECT 126.59 414.18 127.34 414.34 ;
      RECT 121.24 414.1 126.75 414.26 ;
      RECT 121.24 415.06 122.02 415.25 ;
      RECT 121.24 415.06 126.75 415.22 ;
      RECT 126.59 414.98 127.34 415.14 ;
      RECT 126.59 417.58 127.34 417.74 ;
      RECT 121.24 417.5 126.75 417.66 ;
      RECT 121.24 417.47 122.02 417.66 ;
      RECT 121.24 418.46 126.75 418.62 ;
      RECT 126.59 418.38 127.34 418.54 ;
      RECT 126.59 420.98 127.34 421.14 ;
      RECT 121.24 420.9 126.75 421.06 ;
      RECT 121.24 421.86 122.02 422.05 ;
      RECT 121.24 421.86 126.75 422.02 ;
      RECT 126.59 421.78 127.34 421.94 ;
      RECT 126.59 424.38 127.34 424.54 ;
      RECT 121.24 424.3 126.75 424.46 ;
      RECT 121.24 424.27 122.02 424.46 ;
      RECT 121.24 425.26 126.75 425.42 ;
      RECT 126.59 425.18 127.34 425.34 ;
      RECT 126.59 427.78 127.34 427.94 ;
      RECT 121.24 427.7 126.75 427.86 ;
      RECT 121.24 428.66 122.02 428.85 ;
      RECT 121.24 428.66 126.75 428.82 ;
      RECT 126.59 428.58 127.34 428.74 ;
      RECT 126.59 431.18 127.34 431.34 ;
      RECT 121.24 431.1 126.75 431.26 ;
      RECT 121.24 431.07 122.02 431.26 ;
      RECT 121.24 432.06 126.75 432.22 ;
      RECT 126.59 431.98 127.34 432.14 ;
      RECT 126.59 434.58 127.34 434.74 ;
      RECT 121.24 434.5 126.75 434.66 ;
      RECT 121.24 435.46 122.02 435.65 ;
      RECT 121.24 435.46 126.75 435.62 ;
      RECT 126.59 435.38 127.34 435.54 ;
      RECT 126.59 437.98 127.34 438.14 ;
      RECT 121.24 437.9 126.75 438.06 ;
      RECT 121.24 437.87 122.02 438.06 ;
      RECT 121.24 438.86 126.75 439.02 ;
      RECT 126.59 438.78 127.34 438.94 ;
      RECT 126.59 441.38 127.34 441.54 ;
      RECT 121.24 441.3 126.75 441.46 ;
      RECT 121.24 442.26 122.02 442.45 ;
      RECT 121.24 442.26 126.75 442.42 ;
      RECT 126.59 442.18 127.34 442.34 ;
      RECT 126.59 444.78 127.34 444.94 ;
      RECT 121.24 444.7 126.75 444.86 ;
      RECT 121.24 444.67 122.02 444.86 ;
      RECT 121.24 445.66 126.75 445.82 ;
      RECT 126.59 445.58 127.34 445.74 ;
      RECT 126.59 448.18 127.34 448.34 ;
      RECT 121.24 448.1 126.75 448.26 ;
      RECT 121.24 449.06 122.02 449.25 ;
      RECT 121.24 449.06 126.75 449.22 ;
      RECT 126.59 448.98 127.34 449.14 ;
      RECT 126.59 451.58 127.34 451.74 ;
      RECT 121.24 451.5 126.75 451.66 ;
      RECT 121.24 451.47 122.02 451.66 ;
      RECT 121.24 452.46 126.75 452.62 ;
      RECT 126.59 452.38 127.34 452.54 ;
      RECT 126.59 454.98 127.34 455.14 ;
      RECT 121.24 454.9 126.75 455.06 ;
      RECT 121.24 455.86 122.02 456.05 ;
      RECT 121.24 455.86 126.75 456.02 ;
      RECT 126.59 455.78 127.34 455.94 ;
      RECT 126.59 458.38 127.34 458.54 ;
      RECT 121.24 458.3 126.75 458.46 ;
      RECT 121.24 458.27 122.02 458.46 ;
      RECT 121.24 459.26 126.75 459.42 ;
      RECT 126.59 459.18 127.34 459.34 ;
      RECT 126.59 461.78 127.34 461.94 ;
      RECT 121.24 461.7 126.75 461.86 ;
      RECT 121.24 462.66 122.02 462.85 ;
      RECT 121.24 462.66 126.75 462.82 ;
      RECT 126.59 462.58 127.34 462.74 ;
      RECT 126.59 465.18 127.34 465.34 ;
      RECT 121.24 465.1 126.75 465.26 ;
      RECT 121.24 465.07 122.02 465.26 ;
      RECT 121.24 466.06 126.75 466.22 ;
      RECT 126.59 465.98 127.34 466.14 ;
      RECT 126.59 468.58 127.34 468.74 ;
      RECT 121.24 468.5 126.75 468.66 ;
      RECT 121.24 469.46 122.02 469.65 ;
      RECT 121.24 469.46 126.75 469.62 ;
      RECT 126.59 469.38 127.34 469.54 ;
      RECT 126.59 471.98 127.34 472.14 ;
      RECT 121.24 471.9 126.75 472.06 ;
      RECT 121.24 471.87 122.02 472.06 ;
      RECT 121.24 472.86 126.75 473.02 ;
      RECT 126.59 472.78 127.34 472.94 ;
      RECT 126.59 475.38 127.34 475.54 ;
      RECT 121.24 475.3 126.75 475.46 ;
      RECT 121.24 476.26 122.02 476.45 ;
      RECT 121.24 476.26 126.75 476.42 ;
      RECT 126.59 476.18 127.34 476.34 ;
      RECT 126.59 478.78 127.34 478.94 ;
      RECT 121.24 478.7 126.75 478.86 ;
      RECT 121.24 478.67 122.02 478.86 ;
      RECT 121.24 479.66 126.75 479.82 ;
      RECT 126.59 479.58 127.34 479.74 ;
      RECT 126.59 482.18 127.34 482.34 ;
      RECT 121.24 482.1 126.75 482.26 ;
      RECT 121.24 483.06 122.02 483.25 ;
      RECT 121.24 483.06 126.75 483.22 ;
      RECT 126.59 482.98 127.34 483.14 ;
      RECT 126.59 485.58 127.34 485.74 ;
      RECT 121.24 485.5 126.75 485.66 ;
      RECT 121.24 485.47 122.02 485.66 ;
      RECT 121.24 486.46 126.75 486.62 ;
      RECT 126.59 486.38 127.34 486.54 ;
      RECT 126.59 488.98 127.34 489.14 ;
      RECT 121.24 488.9 126.75 489.06 ;
      RECT 121.24 489.86 122.02 490.05 ;
      RECT 121.24 489.86 126.75 490.02 ;
      RECT 126.59 489.78 127.34 489.94 ;
      RECT 126.59 492.38 127.34 492.54 ;
      RECT 121.24 492.3 126.75 492.46 ;
      RECT 121.24 492.27 122.02 492.46 ;
      RECT 121.24 493.26 126.75 493.42 ;
      RECT 126.59 493.18 127.34 493.34 ;
      RECT 126.59 495.78 127.34 495.94 ;
      RECT 121.24 495.7 126.75 495.86 ;
      RECT 121.24 496.66 122.02 496.85 ;
      RECT 121.24 496.66 126.75 496.82 ;
      RECT 126.59 496.58 127.34 496.74 ;
      RECT 126.59 499.18 127.34 499.34 ;
      RECT 121.24 499.1 126.75 499.26 ;
      RECT 121.24 499.07 122.02 499.26 ;
      RECT 121.24 500.06 126.75 500.22 ;
      RECT 126.59 499.98 127.34 500.14 ;
      RECT 126.59 502.58 127.34 502.74 ;
      RECT 121.24 502.5 126.75 502.66 ;
      RECT 121.24 503.46 122.02 503.65 ;
      RECT 121.24 503.46 126.75 503.62 ;
      RECT 126.59 503.38 127.34 503.54 ;
      RECT 126.95 41.08 127.11 45.17 ;
      RECT 126.95 41.08 127.27 41.24 ;
      RECT 126.18 505.54 126.46 506.73 ;
      RECT 125.59 505.54 126.86 505.82 ;
      RECT 126.13 17.6 126.29 23.81 ;
      RECT 125.65 22.38 126.77 22.54 ;
      RECT 126.13 58.24 126.29 64 ;
      RECT 125.65 59.51 126.77 59.67 ;
      RECT 126.55 27.37 126.71 31.49 ;
      RECT 125.71 27.37 125.87 31.49 ;
      RECT 125.71 27.37 126.71 27.53 ;
      RECT 126.13 24.64 126.29 27.53 ;
      RECT 126.13 54.16 126.29 57.42 ;
      RECT 125.71 54.16 126.71 54.88 ;
      RECT 126.55 50.8 126.71 54.88 ;
      RECT 125.71 50.8 125.87 54.88 ;
      RECT 88.11 67.8 126.04 69.03 ;
      RECT 87.75 67.8 126.04 68.69 ;
      RECT 123.97 55.09 125.23 55.25 ;
      RECT 125.07 49.77 125.23 55.25 ;
      RECT 125.07 49.77 125.95 49.93 ;
      RECT 125.79 32.48 125.95 49.93 ;
      RECT 125.13 45.9 125.95 46.06 ;
      RECT 125.13 36.23 125.95 36.39 ;
      RECT 125.07 32.48 125.95 32.64 ;
      RECT 125.07 27.04 125.23 32.64 ;
      RECT 123.97 27.04 125.23 27.2 ;
      RECT 124.86 505.73 125.1 506.76 ;
      RECT 124.86 506.24 125.93 506.51 ;
      RECT 124.64 505.73 125.1 505.96 ;
      RECT 123.87 26.46 125.89 26.62 ;
      RECT 125.73 25.35 125.89 26.62 ;
      RECT 125.65 22.91 125.81 25.51 ;
      RECT 125.65 56.46 125.81 59.14 ;
      RECT 125.73 55.49 125.89 56.62 ;
      RECT 123.87 55.49 125.89 55.65 ;
      RECT 125.33 25.79 125.57 26.07 ;
      RECT 125.33 21.94 125.49 26.07 ;
      RECT 125.33 21.94 125.61 22.18 ;
      RECT 125.39 15.28 125.55 22.18 ;
      RECT 124.43 15.28 124.59 20.88 ;
      RECT 123.47 15.28 123.63 20.88 ;
      RECT 123.47 17.14 125.55 17.3 ;
      RECT 125.39 59.87 125.55 66.77 ;
      RECT 124.43 61.17 124.59 66.77 ;
      RECT 123.47 61.17 123.63 66.77 ;
      RECT 123.47 64.75 125.55 64.91 ;
      RECT 125.33 59.87 125.61 60.11 ;
      RECT 125.33 56.02 125.49 60.11 ;
      RECT 125.33 56.02 125.57 56.3 ;
      RECT 123.47 35.91 125.55 36.07 ;
      RECT 125.39 32.85 125.55 36.07 ;
      RECT 124.43 27.43 124.59 36.07 ;
      RECT 123.47 32.85 123.63 36.07 ;
      RECT 123.53 27.43 124.59 27.59 ;
      RECT 123.53 23.41 123.69 27.59 ;
      RECT 123.53 26.14 124.69 26.3 ;
      RECT 124.53 25.01 124.69 26.3 ;
      RECT 123.53 25 123.73 26.3 ;
      RECT 124.53 21.38 124.69 23.81 ;
      RECT 123.57 21.38 123.73 23.55 ;
      RECT 123.57 21.38 124.69 21.54 ;
      RECT 123.57 60.51 124.69 60.67 ;
      RECT 124.53 58.24 124.69 60.67 ;
      RECT 123.57 58.5 123.73 60.67 ;
      RECT 123.53 55.81 123.69 58.64 ;
      RECT 124.53 55.81 124.69 57.09 ;
      RECT 123.51 55.81 123.73 57.09 ;
      RECT 123.51 55.81 124.69 55.97 ;
      RECT 123.51 54.64 123.67 57.09 ;
      RECT 123.51 54.64 124.59 54.8 ;
      RECT 124.43 46.22 124.59 54.8 ;
      RECT 125.39 46.22 125.55 49.44 ;
      RECT 123.47 46.22 123.63 49.44 ;
      RECT 123.47 46.22 125.55 46.38 ;
      RECT 125.31 41.08 125.47 45.17 ;
      RECT 125.15 41.08 125.47 41.24 ;
      RECT 125.26 505.4 125.42 506.06 ;
      RECT 123.86 505.4 125.42 505.56 ;
      RECT 121.88 505.4 122.74 505.56 ;
      RECT 122.58 505.22 122.74 505.56 ;
      RECT 123.86 505.22 124.02 505.56 ;
      RECT 122.58 505.22 124.02 505.38 ;
      RECT 125.01 21.06 125.17 26.28 ;
      RECT 124.05 24.37 124.21 25.98 ;
      RECT 123.85 24.37 125.17 24.53 ;
      RECT 123.85 23.67 124.01 24.53 ;
      RECT 123.85 23.67 124.21 23.83 ;
      RECT 124.05 21.7 124.21 23.83 ;
      RECT 123.35 21.06 125.23 21.22 ;
      RECT 123.35 60.83 125.23 60.99 ;
      RECT 125.01 55.81 125.17 60.99 ;
      RECT 124.05 58.22 124.21 60.35 ;
      RECT 123.85 58.22 124.21 58.38 ;
      RECT 123.85 57.25 124.01 58.38 ;
      RECT 123.85 57.25 125.17 57.41 ;
      RECT 124.05 56.13 124.21 57.41 ;
      RECT 124.91 32.85 125.07 35.75 ;
      RECT 124.75 31.09 124.91 33.01 ;
      RECT 124.75 49.44 124.91 51.3 ;
      RECT 124.91 46.54 125.07 49.6 ;
      RECT 124.83 38.57 124.99 45.17 ;
      RECT 124.53 38.57 124.99 38.73 ;
      RECT 124.53 36.23 124.69 38.73 ;
      RECT 124.17 36.23 124.85 36.39 ;
      RECT 124.05 45.9 124.85 46.06 ;
      RECT 124.05 44.89 124.21 46.06 ;
      RECT 124.03 38.57 124.19 45.17 ;
      RECT 124.08 70.38 124.7 70.54 ;
      RECT 124.08 69.85 124.24 70.54 ;
      RECT 121.74 69.96 123.06 70.12 ;
      RECT 122.88 69.85 124.24 70.02 ;
      RECT 122.88 75.9 124.24 76.07 ;
      RECT 124.08 75.38 124.24 76.07 ;
      RECT 121.74 75.8 123.06 75.96 ;
      RECT 124.08 75.38 124.7 75.54 ;
      RECT 124.08 77.18 124.7 77.34 ;
      RECT 124.08 76.65 124.24 77.34 ;
      RECT 121.74 76.76 123.06 76.92 ;
      RECT 122.88 76.65 124.24 76.82 ;
      RECT 122.88 82.7 124.24 82.87 ;
      RECT 124.08 82.18 124.24 82.87 ;
      RECT 121.74 82.6 123.06 82.76 ;
      RECT 124.08 82.18 124.7 82.34 ;
      RECT 124.08 83.98 124.7 84.14 ;
      RECT 124.08 83.45 124.24 84.14 ;
      RECT 121.74 83.56 123.06 83.72 ;
      RECT 122.88 83.45 124.24 83.62 ;
      RECT 122.88 89.5 124.24 89.67 ;
      RECT 124.08 88.98 124.24 89.67 ;
      RECT 121.74 89.4 123.06 89.56 ;
      RECT 124.08 88.98 124.7 89.14 ;
      RECT 124.08 90.78 124.7 90.94 ;
      RECT 124.08 90.25 124.24 90.94 ;
      RECT 121.74 90.36 123.06 90.52 ;
      RECT 122.88 90.25 124.24 90.42 ;
      RECT 122.88 96.3 124.24 96.47 ;
      RECT 124.08 95.78 124.24 96.47 ;
      RECT 121.74 96.2 123.06 96.36 ;
      RECT 124.08 95.78 124.7 95.94 ;
      RECT 124.08 97.58 124.7 97.74 ;
      RECT 124.08 97.05 124.24 97.74 ;
      RECT 121.74 97.16 123.06 97.32 ;
      RECT 122.88 97.05 124.24 97.22 ;
      RECT 122.88 103.1 124.24 103.27 ;
      RECT 124.08 102.58 124.24 103.27 ;
      RECT 121.74 103 123.06 103.16 ;
      RECT 124.08 102.58 124.7 102.74 ;
      RECT 124.08 104.38 124.7 104.54 ;
      RECT 124.08 103.85 124.24 104.54 ;
      RECT 121.74 103.96 123.06 104.12 ;
      RECT 122.88 103.85 124.24 104.02 ;
      RECT 122.88 109.9 124.24 110.07 ;
      RECT 124.08 109.38 124.24 110.07 ;
      RECT 121.74 109.8 123.06 109.96 ;
      RECT 124.08 109.38 124.7 109.54 ;
      RECT 124.08 111.18 124.7 111.34 ;
      RECT 124.08 110.65 124.24 111.34 ;
      RECT 121.74 110.76 123.06 110.92 ;
      RECT 122.88 110.65 124.24 110.82 ;
      RECT 122.88 116.7 124.24 116.87 ;
      RECT 124.08 116.18 124.24 116.87 ;
      RECT 121.74 116.6 123.06 116.76 ;
      RECT 124.08 116.18 124.7 116.34 ;
      RECT 124.08 117.98 124.7 118.14 ;
      RECT 124.08 117.45 124.24 118.14 ;
      RECT 121.74 117.56 123.06 117.72 ;
      RECT 122.88 117.45 124.24 117.62 ;
      RECT 122.88 123.5 124.24 123.67 ;
      RECT 124.08 122.98 124.24 123.67 ;
      RECT 121.74 123.4 123.06 123.56 ;
      RECT 124.08 122.98 124.7 123.14 ;
      RECT 124.08 124.78 124.7 124.94 ;
      RECT 124.08 124.25 124.24 124.94 ;
      RECT 121.74 124.36 123.06 124.52 ;
      RECT 122.88 124.25 124.24 124.42 ;
      RECT 122.88 130.3 124.24 130.47 ;
      RECT 124.08 129.78 124.24 130.47 ;
      RECT 121.74 130.2 123.06 130.36 ;
      RECT 124.08 129.78 124.7 129.94 ;
      RECT 124.08 131.58 124.7 131.74 ;
      RECT 124.08 131.05 124.24 131.74 ;
      RECT 121.74 131.16 123.06 131.32 ;
      RECT 122.88 131.05 124.24 131.22 ;
      RECT 122.88 137.1 124.24 137.27 ;
      RECT 124.08 136.58 124.24 137.27 ;
      RECT 121.74 137 123.06 137.16 ;
      RECT 124.08 136.58 124.7 136.74 ;
      RECT 124.08 138.38 124.7 138.54 ;
      RECT 124.08 137.85 124.24 138.54 ;
      RECT 121.74 137.96 123.06 138.12 ;
      RECT 122.88 137.85 124.24 138.02 ;
      RECT 122.88 143.9 124.24 144.07 ;
      RECT 124.08 143.38 124.24 144.07 ;
      RECT 121.74 143.8 123.06 143.96 ;
      RECT 124.08 143.38 124.7 143.54 ;
      RECT 124.08 145.18 124.7 145.34 ;
      RECT 124.08 144.65 124.24 145.34 ;
      RECT 121.74 144.76 123.06 144.92 ;
      RECT 122.88 144.65 124.24 144.82 ;
      RECT 122.88 150.7 124.24 150.87 ;
      RECT 124.08 150.18 124.24 150.87 ;
      RECT 121.74 150.6 123.06 150.76 ;
      RECT 124.08 150.18 124.7 150.34 ;
      RECT 124.08 151.98 124.7 152.14 ;
      RECT 124.08 151.45 124.24 152.14 ;
      RECT 121.74 151.56 123.06 151.72 ;
      RECT 122.88 151.45 124.24 151.62 ;
      RECT 122.88 157.5 124.24 157.67 ;
      RECT 124.08 156.98 124.24 157.67 ;
      RECT 121.74 157.4 123.06 157.56 ;
      RECT 124.08 156.98 124.7 157.14 ;
      RECT 124.08 158.78 124.7 158.94 ;
      RECT 124.08 158.25 124.24 158.94 ;
      RECT 121.74 158.36 123.06 158.52 ;
      RECT 122.88 158.25 124.24 158.42 ;
      RECT 122.88 164.3 124.24 164.47 ;
      RECT 124.08 163.78 124.24 164.47 ;
      RECT 121.74 164.2 123.06 164.36 ;
      RECT 124.08 163.78 124.7 163.94 ;
      RECT 124.08 165.58 124.7 165.74 ;
      RECT 124.08 165.05 124.24 165.74 ;
      RECT 121.74 165.16 123.06 165.32 ;
      RECT 122.88 165.05 124.24 165.22 ;
      RECT 122.88 171.1 124.24 171.27 ;
      RECT 124.08 170.58 124.24 171.27 ;
      RECT 121.74 171 123.06 171.16 ;
      RECT 124.08 170.58 124.7 170.74 ;
      RECT 124.08 172.38 124.7 172.54 ;
      RECT 124.08 171.85 124.24 172.54 ;
      RECT 121.74 171.96 123.06 172.12 ;
      RECT 122.88 171.85 124.24 172.02 ;
      RECT 122.88 177.9 124.24 178.07 ;
      RECT 124.08 177.38 124.24 178.07 ;
      RECT 121.74 177.8 123.06 177.96 ;
      RECT 124.08 177.38 124.7 177.54 ;
      RECT 124.08 179.18 124.7 179.34 ;
      RECT 124.08 178.65 124.24 179.34 ;
      RECT 121.74 178.76 123.06 178.92 ;
      RECT 122.88 178.65 124.24 178.82 ;
      RECT 122.88 184.7 124.24 184.87 ;
      RECT 124.08 184.18 124.24 184.87 ;
      RECT 121.74 184.6 123.06 184.76 ;
      RECT 124.08 184.18 124.7 184.34 ;
      RECT 124.08 185.98 124.7 186.14 ;
      RECT 124.08 185.45 124.24 186.14 ;
      RECT 121.74 185.56 123.06 185.72 ;
      RECT 122.88 185.45 124.24 185.62 ;
      RECT 122.88 191.5 124.24 191.67 ;
      RECT 124.08 190.98 124.24 191.67 ;
      RECT 121.74 191.4 123.06 191.56 ;
      RECT 124.08 190.98 124.7 191.14 ;
      RECT 124.08 192.78 124.7 192.94 ;
      RECT 124.08 192.25 124.24 192.94 ;
      RECT 121.74 192.36 123.06 192.52 ;
      RECT 122.88 192.25 124.24 192.42 ;
      RECT 122.88 198.3 124.24 198.47 ;
      RECT 124.08 197.78 124.24 198.47 ;
      RECT 121.74 198.2 123.06 198.36 ;
      RECT 124.08 197.78 124.7 197.94 ;
      RECT 124.08 199.58 124.7 199.74 ;
      RECT 124.08 199.05 124.24 199.74 ;
      RECT 121.74 199.16 123.06 199.32 ;
      RECT 122.88 199.05 124.24 199.22 ;
      RECT 122.88 205.1 124.24 205.27 ;
      RECT 124.08 204.58 124.24 205.27 ;
      RECT 121.74 205 123.06 205.16 ;
      RECT 124.08 204.58 124.7 204.74 ;
      RECT 124.08 206.38 124.7 206.54 ;
      RECT 124.08 205.85 124.24 206.54 ;
      RECT 121.74 205.96 123.06 206.12 ;
      RECT 122.88 205.85 124.24 206.02 ;
      RECT 122.88 211.9 124.24 212.07 ;
      RECT 124.08 211.38 124.24 212.07 ;
      RECT 121.74 211.8 123.06 211.96 ;
      RECT 124.08 211.38 124.7 211.54 ;
      RECT 124.08 213.18 124.7 213.34 ;
      RECT 124.08 212.65 124.24 213.34 ;
      RECT 121.74 212.76 123.06 212.92 ;
      RECT 122.88 212.65 124.24 212.82 ;
      RECT 122.88 218.7 124.24 218.87 ;
      RECT 124.08 218.18 124.24 218.87 ;
      RECT 121.74 218.6 123.06 218.76 ;
      RECT 124.08 218.18 124.7 218.34 ;
      RECT 124.08 219.98 124.7 220.14 ;
      RECT 124.08 219.45 124.24 220.14 ;
      RECT 121.74 219.56 123.06 219.72 ;
      RECT 122.88 219.45 124.24 219.62 ;
      RECT 122.88 225.5 124.24 225.67 ;
      RECT 124.08 224.98 124.24 225.67 ;
      RECT 121.74 225.4 123.06 225.56 ;
      RECT 124.08 224.98 124.7 225.14 ;
      RECT 124.08 226.78 124.7 226.94 ;
      RECT 124.08 226.25 124.24 226.94 ;
      RECT 121.74 226.36 123.06 226.52 ;
      RECT 122.88 226.25 124.24 226.42 ;
      RECT 122.88 232.3 124.24 232.47 ;
      RECT 124.08 231.78 124.24 232.47 ;
      RECT 121.74 232.2 123.06 232.36 ;
      RECT 124.08 231.78 124.7 231.94 ;
      RECT 124.08 233.58 124.7 233.74 ;
      RECT 124.08 233.05 124.24 233.74 ;
      RECT 121.74 233.16 123.06 233.32 ;
      RECT 122.88 233.05 124.24 233.22 ;
      RECT 122.88 239.1 124.24 239.27 ;
      RECT 124.08 238.58 124.24 239.27 ;
      RECT 121.74 239 123.06 239.16 ;
      RECT 124.08 238.58 124.7 238.74 ;
      RECT 124.08 240.38 124.7 240.54 ;
      RECT 124.08 239.85 124.24 240.54 ;
      RECT 121.74 239.96 123.06 240.12 ;
      RECT 122.88 239.85 124.24 240.02 ;
      RECT 122.88 245.9 124.24 246.07 ;
      RECT 124.08 245.38 124.24 246.07 ;
      RECT 121.74 245.8 123.06 245.96 ;
      RECT 124.08 245.38 124.7 245.54 ;
      RECT 124.08 247.18 124.7 247.34 ;
      RECT 124.08 246.65 124.24 247.34 ;
      RECT 121.74 246.76 123.06 246.92 ;
      RECT 122.88 246.65 124.24 246.82 ;
      RECT 122.88 252.7 124.24 252.87 ;
      RECT 124.08 252.18 124.24 252.87 ;
      RECT 121.74 252.6 123.06 252.76 ;
      RECT 124.08 252.18 124.7 252.34 ;
      RECT 124.08 253.98 124.7 254.14 ;
      RECT 124.08 253.45 124.24 254.14 ;
      RECT 121.74 253.56 123.06 253.72 ;
      RECT 122.88 253.45 124.24 253.62 ;
      RECT 122.88 259.5 124.24 259.67 ;
      RECT 124.08 258.98 124.24 259.67 ;
      RECT 121.74 259.4 123.06 259.56 ;
      RECT 124.08 258.98 124.7 259.14 ;
      RECT 124.08 260.78 124.7 260.94 ;
      RECT 124.08 260.25 124.24 260.94 ;
      RECT 121.74 260.36 123.06 260.52 ;
      RECT 122.88 260.25 124.24 260.42 ;
      RECT 122.88 266.3 124.24 266.47 ;
      RECT 124.08 265.78 124.24 266.47 ;
      RECT 121.74 266.2 123.06 266.36 ;
      RECT 124.08 265.78 124.7 265.94 ;
      RECT 124.08 267.58 124.7 267.74 ;
      RECT 124.08 267.05 124.24 267.74 ;
      RECT 121.74 267.16 123.06 267.32 ;
      RECT 122.88 267.05 124.24 267.22 ;
      RECT 122.88 273.1 124.24 273.27 ;
      RECT 124.08 272.58 124.24 273.27 ;
      RECT 121.74 273 123.06 273.16 ;
      RECT 124.08 272.58 124.7 272.74 ;
      RECT 124.08 274.38 124.7 274.54 ;
      RECT 124.08 273.85 124.24 274.54 ;
      RECT 121.74 273.96 123.06 274.12 ;
      RECT 122.88 273.85 124.24 274.02 ;
      RECT 122.88 279.9 124.24 280.07 ;
      RECT 124.08 279.38 124.24 280.07 ;
      RECT 121.74 279.8 123.06 279.96 ;
      RECT 124.08 279.38 124.7 279.54 ;
      RECT 124.08 281.18 124.7 281.34 ;
      RECT 124.08 280.65 124.24 281.34 ;
      RECT 121.74 280.76 123.06 280.92 ;
      RECT 122.88 280.65 124.24 280.82 ;
      RECT 122.88 286.7 124.24 286.87 ;
      RECT 124.08 286.18 124.24 286.87 ;
      RECT 121.74 286.6 123.06 286.76 ;
      RECT 124.08 286.18 124.7 286.34 ;
      RECT 124.08 287.98 124.7 288.14 ;
      RECT 124.08 287.45 124.24 288.14 ;
      RECT 121.74 287.56 123.06 287.72 ;
      RECT 122.88 287.45 124.24 287.62 ;
      RECT 122.88 293.5 124.24 293.67 ;
      RECT 124.08 292.98 124.24 293.67 ;
      RECT 121.74 293.4 123.06 293.56 ;
      RECT 124.08 292.98 124.7 293.14 ;
      RECT 124.08 294.78 124.7 294.94 ;
      RECT 124.08 294.25 124.24 294.94 ;
      RECT 121.74 294.36 123.06 294.52 ;
      RECT 122.88 294.25 124.24 294.42 ;
      RECT 122.88 300.3 124.24 300.47 ;
      RECT 124.08 299.78 124.24 300.47 ;
      RECT 121.74 300.2 123.06 300.36 ;
      RECT 124.08 299.78 124.7 299.94 ;
      RECT 124.08 301.58 124.7 301.74 ;
      RECT 124.08 301.05 124.24 301.74 ;
      RECT 121.74 301.16 123.06 301.32 ;
      RECT 122.88 301.05 124.24 301.22 ;
      RECT 122.88 307.1 124.24 307.27 ;
      RECT 124.08 306.58 124.24 307.27 ;
      RECT 121.74 307 123.06 307.16 ;
      RECT 124.08 306.58 124.7 306.74 ;
      RECT 124.08 308.38 124.7 308.54 ;
      RECT 124.08 307.85 124.24 308.54 ;
      RECT 121.74 307.96 123.06 308.12 ;
      RECT 122.88 307.85 124.24 308.02 ;
      RECT 122.88 313.9 124.24 314.07 ;
      RECT 124.08 313.38 124.24 314.07 ;
      RECT 121.74 313.8 123.06 313.96 ;
      RECT 124.08 313.38 124.7 313.54 ;
      RECT 124.08 315.18 124.7 315.34 ;
      RECT 124.08 314.65 124.24 315.34 ;
      RECT 121.74 314.76 123.06 314.92 ;
      RECT 122.88 314.65 124.24 314.82 ;
      RECT 122.88 320.7 124.24 320.87 ;
      RECT 124.08 320.18 124.24 320.87 ;
      RECT 121.74 320.6 123.06 320.76 ;
      RECT 124.08 320.18 124.7 320.34 ;
      RECT 124.08 321.98 124.7 322.14 ;
      RECT 124.08 321.45 124.24 322.14 ;
      RECT 121.74 321.56 123.06 321.72 ;
      RECT 122.88 321.45 124.24 321.62 ;
      RECT 122.88 327.5 124.24 327.67 ;
      RECT 124.08 326.98 124.24 327.67 ;
      RECT 121.74 327.4 123.06 327.56 ;
      RECT 124.08 326.98 124.7 327.14 ;
      RECT 124.08 328.78 124.7 328.94 ;
      RECT 124.08 328.25 124.24 328.94 ;
      RECT 121.74 328.36 123.06 328.52 ;
      RECT 122.88 328.25 124.24 328.42 ;
      RECT 122.88 334.3 124.24 334.47 ;
      RECT 124.08 333.78 124.24 334.47 ;
      RECT 121.74 334.2 123.06 334.36 ;
      RECT 124.08 333.78 124.7 333.94 ;
      RECT 124.08 335.58 124.7 335.74 ;
      RECT 124.08 335.05 124.24 335.74 ;
      RECT 121.74 335.16 123.06 335.32 ;
      RECT 122.88 335.05 124.24 335.22 ;
      RECT 122.88 341.1 124.24 341.27 ;
      RECT 124.08 340.58 124.24 341.27 ;
      RECT 121.74 341 123.06 341.16 ;
      RECT 124.08 340.58 124.7 340.74 ;
      RECT 124.08 342.38 124.7 342.54 ;
      RECT 124.08 341.85 124.24 342.54 ;
      RECT 121.74 341.96 123.06 342.12 ;
      RECT 122.88 341.85 124.24 342.02 ;
      RECT 122.88 347.9 124.24 348.07 ;
      RECT 124.08 347.38 124.24 348.07 ;
      RECT 121.74 347.8 123.06 347.96 ;
      RECT 124.08 347.38 124.7 347.54 ;
      RECT 124.08 349.18 124.7 349.34 ;
      RECT 124.08 348.65 124.24 349.34 ;
      RECT 121.74 348.76 123.06 348.92 ;
      RECT 122.88 348.65 124.24 348.82 ;
      RECT 122.88 354.7 124.24 354.87 ;
      RECT 124.08 354.18 124.24 354.87 ;
      RECT 121.74 354.6 123.06 354.76 ;
      RECT 124.08 354.18 124.7 354.34 ;
      RECT 124.08 355.98 124.7 356.14 ;
      RECT 124.08 355.45 124.24 356.14 ;
      RECT 121.74 355.56 123.06 355.72 ;
      RECT 122.88 355.45 124.24 355.62 ;
      RECT 122.88 361.5 124.24 361.67 ;
      RECT 124.08 360.98 124.24 361.67 ;
      RECT 121.74 361.4 123.06 361.56 ;
      RECT 124.08 360.98 124.7 361.14 ;
      RECT 124.08 362.78 124.7 362.94 ;
      RECT 124.08 362.25 124.24 362.94 ;
      RECT 121.74 362.36 123.06 362.52 ;
      RECT 122.88 362.25 124.24 362.42 ;
      RECT 122.88 368.3 124.24 368.47 ;
      RECT 124.08 367.78 124.24 368.47 ;
      RECT 121.74 368.2 123.06 368.36 ;
      RECT 124.08 367.78 124.7 367.94 ;
      RECT 124.08 369.58 124.7 369.74 ;
      RECT 124.08 369.05 124.24 369.74 ;
      RECT 121.74 369.16 123.06 369.32 ;
      RECT 122.88 369.05 124.24 369.22 ;
      RECT 122.88 375.1 124.24 375.27 ;
      RECT 124.08 374.58 124.24 375.27 ;
      RECT 121.74 375 123.06 375.16 ;
      RECT 124.08 374.58 124.7 374.74 ;
      RECT 124.08 376.38 124.7 376.54 ;
      RECT 124.08 375.85 124.24 376.54 ;
      RECT 121.74 375.96 123.06 376.12 ;
      RECT 122.88 375.85 124.24 376.02 ;
      RECT 122.88 381.9 124.24 382.07 ;
      RECT 124.08 381.38 124.24 382.07 ;
      RECT 121.74 381.8 123.06 381.96 ;
      RECT 124.08 381.38 124.7 381.54 ;
      RECT 124.08 383.18 124.7 383.34 ;
      RECT 124.08 382.65 124.24 383.34 ;
      RECT 121.74 382.76 123.06 382.92 ;
      RECT 122.88 382.65 124.24 382.82 ;
      RECT 122.88 388.7 124.24 388.87 ;
      RECT 124.08 388.18 124.24 388.87 ;
      RECT 121.74 388.6 123.06 388.76 ;
      RECT 124.08 388.18 124.7 388.34 ;
      RECT 124.08 389.98 124.7 390.14 ;
      RECT 124.08 389.45 124.24 390.14 ;
      RECT 121.74 389.56 123.06 389.72 ;
      RECT 122.88 389.45 124.24 389.62 ;
      RECT 122.88 395.5 124.24 395.67 ;
      RECT 124.08 394.98 124.24 395.67 ;
      RECT 121.74 395.4 123.06 395.56 ;
      RECT 124.08 394.98 124.7 395.14 ;
      RECT 124.08 396.78 124.7 396.94 ;
      RECT 124.08 396.25 124.24 396.94 ;
      RECT 121.74 396.36 123.06 396.52 ;
      RECT 122.88 396.25 124.24 396.42 ;
      RECT 122.88 402.3 124.24 402.47 ;
      RECT 124.08 401.78 124.24 402.47 ;
      RECT 121.74 402.2 123.06 402.36 ;
      RECT 124.08 401.78 124.7 401.94 ;
      RECT 124.08 403.58 124.7 403.74 ;
      RECT 124.08 403.05 124.24 403.74 ;
      RECT 121.74 403.16 123.06 403.32 ;
      RECT 122.88 403.05 124.24 403.22 ;
      RECT 122.88 409.1 124.24 409.27 ;
      RECT 124.08 408.58 124.24 409.27 ;
      RECT 121.74 409 123.06 409.16 ;
      RECT 124.08 408.58 124.7 408.74 ;
      RECT 124.08 410.38 124.7 410.54 ;
      RECT 124.08 409.85 124.24 410.54 ;
      RECT 121.74 409.96 123.06 410.12 ;
      RECT 122.88 409.85 124.24 410.02 ;
      RECT 122.88 415.9 124.24 416.07 ;
      RECT 124.08 415.38 124.24 416.07 ;
      RECT 121.74 415.8 123.06 415.96 ;
      RECT 124.08 415.38 124.7 415.54 ;
      RECT 124.08 417.18 124.7 417.34 ;
      RECT 124.08 416.65 124.24 417.34 ;
      RECT 121.74 416.76 123.06 416.92 ;
      RECT 122.88 416.65 124.24 416.82 ;
      RECT 122.88 422.7 124.24 422.87 ;
      RECT 124.08 422.18 124.24 422.87 ;
      RECT 121.74 422.6 123.06 422.76 ;
      RECT 124.08 422.18 124.7 422.34 ;
      RECT 124.08 423.98 124.7 424.14 ;
      RECT 124.08 423.45 124.24 424.14 ;
      RECT 121.74 423.56 123.06 423.72 ;
      RECT 122.88 423.45 124.24 423.62 ;
      RECT 122.88 429.5 124.24 429.67 ;
      RECT 124.08 428.98 124.24 429.67 ;
      RECT 121.74 429.4 123.06 429.56 ;
      RECT 124.08 428.98 124.7 429.14 ;
      RECT 124.08 430.78 124.7 430.94 ;
      RECT 124.08 430.25 124.24 430.94 ;
      RECT 121.74 430.36 123.06 430.52 ;
      RECT 122.88 430.25 124.24 430.42 ;
      RECT 122.88 436.3 124.24 436.47 ;
      RECT 124.08 435.78 124.24 436.47 ;
      RECT 121.74 436.2 123.06 436.36 ;
      RECT 124.08 435.78 124.7 435.94 ;
      RECT 124.08 437.58 124.7 437.74 ;
      RECT 124.08 437.05 124.24 437.74 ;
      RECT 121.74 437.16 123.06 437.32 ;
      RECT 122.88 437.05 124.24 437.22 ;
      RECT 122.88 443.1 124.24 443.27 ;
      RECT 124.08 442.58 124.24 443.27 ;
      RECT 121.74 443 123.06 443.16 ;
      RECT 124.08 442.58 124.7 442.74 ;
      RECT 124.08 444.38 124.7 444.54 ;
      RECT 124.08 443.85 124.24 444.54 ;
      RECT 121.74 443.96 123.06 444.12 ;
      RECT 122.88 443.85 124.24 444.02 ;
      RECT 122.88 449.9 124.24 450.07 ;
      RECT 124.08 449.38 124.24 450.07 ;
      RECT 121.74 449.8 123.06 449.96 ;
      RECT 124.08 449.38 124.7 449.54 ;
      RECT 124.08 451.18 124.7 451.34 ;
      RECT 124.08 450.65 124.24 451.34 ;
      RECT 121.74 450.76 123.06 450.92 ;
      RECT 122.88 450.65 124.24 450.82 ;
      RECT 122.88 456.7 124.24 456.87 ;
      RECT 124.08 456.18 124.24 456.87 ;
      RECT 121.74 456.6 123.06 456.76 ;
      RECT 124.08 456.18 124.7 456.34 ;
      RECT 124.08 457.98 124.7 458.14 ;
      RECT 124.08 457.45 124.24 458.14 ;
      RECT 121.74 457.56 123.06 457.72 ;
      RECT 122.88 457.45 124.24 457.62 ;
      RECT 122.88 463.5 124.24 463.67 ;
      RECT 124.08 462.98 124.24 463.67 ;
      RECT 121.74 463.4 123.06 463.56 ;
      RECT 124.08 462.98 124.7 463.14 ;
      RECT 124.08 464.78 124.7 464.94 ;
      RECT 124.08 464.25 124.24 464.94 ;
      RECT 121.74 464.36 123.06 464.52 ;
      RECT 122.88 464.25 124.24 464.42 ;
      RECT 122.88 470.3 124.24 470.47 ;
      RECT 124.08 469.78 124.24 470.47 ;
      RECT 121.74 470.2 123.06 470.36 ;
      RECT 124.08 469.78 124.7 469.94 ;
      RECT 124.08 471.58 124.7 471.74 ;
      RECT 124.08 471.05 124.24 471.74 ;
      RECT 121.74 471.16 123.06 471.32 ;
      RECT 122.88 471.05 124.24 471.22 ;
      RECT 122.88 477.1 124.24 477.27 ;
      RECT 124.08 476.58 124.24 477.27 ;
      RECT 121.74 477 123.06 477.16 ;
      RECT 124.08 476.58 124.7 476.74 ;
      RECT 124.08 478.38 124.7 478.54 ;
      RECT 124.08 477.85 124.24 478.54 ;
      RECT 121.74 477.96 123.06 478.12 ;
      RECT 122.88 477.85 124.24 478.02 ;
      RECT 122.88 483.9 124.24 484.07 ;
      RECT 124.08 483.38 124.24 484.07 ;
      RECT 121.74 483.8 123.06 483.96 ;
      RECT 124.08 483.38 124.7 483.54 ;
      RECT 124.08 485.18 124.7 485.34 ;
      RECT 124.08 484.65 124.24 485.34 ;
      RECT 121.74 484.76 123.06 484.92 ;
      RECT 122.88 484.65 124.24 484.82 ;
      RECT 122.88 490.7 124.24 490.87 ;
      RECT 124.08 490.18 124.24 490.87 ;
      RECT 121.74 490.6 123.06 490.76 ;
      RECT 124.08 490.18 124.7 490.34 ;
      RECT 124.08 491.98 124.7 492.14 ;
      RECT 124.08 491.45 124.24 492.14 ;
      RECT 121.74 491.56 123.06 491.72 ;
      RECT 122.88 491.45 124.24 491.62 ;
      RECT 122.88 497.5 124.24 497.67 ;
      RECT 124.08 496.98 124.24 497.67 ;
      RECT 121.74 497.4 123.06 497.56 ;
      RECT 124.08 496.98 124.7 497.14 ;
      RECT 124.08 498.78 124.7 498.94 ;
      RECT 124.08 498.25 124.24 498.94 ;
      RECT 121.74 498.36 123.06 498.52 ;
      RECT 122.88 498.25 124.24 498.42 ;
      RECT 122.88 504.3 124.24 504.47 ;
      RECT 124.08 503.78 124.24 504.47 ;
      RECT 121.74 504.2 123.06 504.36 ;
      RECT 124.08 503.78 124.7 503.94 ;
      RECT 121.76 72.5 124.22 72.66 ;
      RECT 124.06 71.98 124.22 72.66 ;
      RECT 121.66 72.4 121.94 72.56 ;
      RECT 124.06 71.98 124.68 72.14 ;
      RECT 124.06 73.78 124.68 73.94 ;
      RECT 124.06 73.26 124.22 73.94 ;
      RECT 121.66 73.36 121.94 73.52 ;
      RECT 121.76 73.26 124.22 73.42 ;
      RECT 121.76 79.3 124.22 79.46 ;
      RECT 124.06 78.78 124.22 79.46 ;
      RECT 121.66 79.2 121.94 79.36 ;
      RECT 124.06 78.78 124.68 78.94 ;
      RECT 124.06 80.58 124.68 80.74 ;
      RECT 124.06 80.06 124.22 80.74 ;
      RECT 121.66 80.16 121.94 80.32 ;
      RECT 121.76 80.06 124.22 80.22 ;
      RECT 121.76 86.1 124.22 86.26 ;
      RECT 124.06 85.58 124.22 86.26 ;
      RECT 121.66 86 121.94 86.16 ;
      RECT 124.06 85.58 124.68 85.74 ;
      RECT 124.06 87.38 124.68 87.54 ;
      RECT 124.06 86.86 124.22 87.54 ;
      RECT 121.66 86.96 121.94 87.12 ;
      RECT 121.76 86.86 124.22 87.02 ;
      RECT 121.76 92.9 124.22 93.06 ;
      RECT 124.06 92.38 124.22 93.06 ;
      RECT 121.66 92.8 121.94 92.96 ;
      RECT 124.06 92.38 124.68 92.54 ;
      RECT 124.06 94.18 124.68 94.34 ;
      RECT 124.06 93.66 124.22 94.34 ;
      RECT 121.66 93.76 121.94 93.92 ;
      RECT 121.76 93.66 124.22 93.82 ;
      RECT 121.76 99.7 124.22 99.86 ;
      RECT 124.06 99.18 124.22 99.86 ;
      RECT 121.66 99.6 121.94 99.76 ;
      RECT 124.06 99.18 124.68 99.34 ;
      RECT 124.06 100.98 124.68 101.14 ;
      RECT 124.06 100.46 124.22 101.14 ;
      RECT 121.66 100.56 121.94 100.72 ;
      RECT 121.76 100.46 124.22 100.62 ;
      RECT 121.76 106.5 124.22 106.66 ;
      RECT 124.06 105.98 124.22 106.66 ;
      RECT 121.66 106.4 121.94 106.56 ;
      RECT 124.06 105.98 124.68 106.14 ;
      RECT 124.06 107.78 124.68 107.94 ;
      RECT 124.06 107.26 124.22 107.94 ;
      RECT 121.66 107.36 121.94 107.52 ;
      RECT 121.76 107.26 124.22 107.42 ;
      RECT 121.76 113.3 124.22 113.46 ;
      RECT 124.06 112.78 124.22 113.46 ;
      RECT 121.66 113.2 121.94 113.36 ;
      RECT 124.06 112.78 124.68 112.94 ;
      RECT 124.06 114.58 124.68 114.74 ;
      RECT 124.06 114.06 124.22 114.74 ;
      RECT 121.66 114.16 121.94 114.32 ;
      RECT 121.76 114.06 124.22 114.22 ;
      RECT 121.76 120.1 124.22 120.26 ;
      RECT 124.06 119.58 124.22 120.26 ;
      RECT 121.66 120 121.94 120.16 ;
      RECT 124.06 119.58 124.68 119.74 ;
      RECT 124.06 121.38 124.68 121.54 ;
      RECT 124.06 120.86 124.22 121.54 ;
      RECT 121.66 120.96 121.94 121.12 ;
      RECT 121.76 120.86 124.22 121.02 ;
      RECT 121.76 126.9 124.22 127.06 ;
      RECT 124.06 126.38 124.22 127.06 ;
      RECT 121.66 126.8 121.94 126.96 ;
      RECT 124.06 126.38 124.68 126.54 ;
      RECT 124.06 128.18 124.68 128.34 ;
      RECT 124.06 127.66 124.22 128.34 ;
      RECT 121.66 127.76 121.94 127.92 ;
      RECT 121.76 127.66 124.22 127.82 ;
      RECT 121.76 133.7 124.22 133.86 ;
      RECT 124.06 133.18 124.22 133.86 ;
      RECT 121.66 133.6 121.94 133.76 ;
      RECT 124.06 133.18 124.68 133.34 ;
      RECT 124.06 134.98 124.68 135.14 ;
      RECT 124.06 134.46 124.22 135.14 ;
      RECT 121.66 134.56 121.94 134.72 ;
      RECT 121.76 134.46 124.22 134.62 ;
      RECT 121.76 140.5 124.22 140.66 ;
      RECT 124.06 139.98 124.22 140.66 ;
      RECT 121.66 140.4 121.94 140.56 ;
      RECT 124.06 139.98 124.68 140.14 ;
      RECT 124.06 141.78 124.68 141.94 ;
      RECT 124.06 141.26 124.22 141.94 ;
      RECT 121.66 141.36 121.94 141.52 ;
      RECT 121.76 141.26 124.22 141.42 ;
      RECT 121.76 147.3 124.22 147.46 ;
      RECT 124.06 146.78 124.22 147.46 ;
      RECT 121.66 147.2 121.94 147.36 ;
      RECT 124.06 146.78 124.68 146.94 ;
      RECT 124.06 148.58 124.68 148.74 ;
      RECT 124.06 148.06 124.22 148.74 ;
      RECT 121.66 148.16 121.94 148.32 ;
      RECT 121.76 148.06 124.22 148.22 ;
      RECT 121.76 154.1 124.22 154.26 ;
      RECT 124.06 153.58 124.22 154.26 ;
      RECT 121.66 154 121.94 154.16 ;
      RECT 124.06 153.58 124.68 153.74 ;
      RECT 124.06 155.38 124.68 155.54 ;
      RECT 124.06 154.86 124.22 155.54 ;
      RECT 121.66 154.96 121.94 155.12 ;
      RECT 121.76 154.86 124.22 155.02 ;
      RECT 121.76 160.9 124.22 161.06 ;
      RECT 124.06 160.38 124.22 161.06 ;
      RECT 121.66 160.8 121.94 160.96 ;
      RECT 124.06 160.38 124.68 160.54 ;
      RECT 124.06 162.18 124.68 162.34 ;
      RECT 124.06 161.66 124.22 162.34 ;
      RECT 121.66 161.76 121.94 161.92 ;
      RECT 121.76 161.66 124.22 161.82 ;
      RECT 121.76 167.7 124.22 167.86 ;
      RECT 124.06 167.18 124.22 167.86 ;
      RECT 121.66 167.6 121.94 167.76 ;
      RECT 124.06 167.18 124.68 167.34 ;
      RECT 124.06 168.98 124.68 169.14 ;
      RECT 124.06 168.46 124.22 169.14 ;
      RECT 121.66 168.56 121.94 168.72 ;
      RECT 121.76 168.46 124.22 168.62 ;
      RECT 121.76 174.5 124.22 174.66 ;
      RECT 124.06 173.98 124.22 174.66 ;
      RECT 121.66 174.4 121.94 174.56 ;
      RECT 124.06 173.98 124.68 174.14 ;
      RECT 124.06 175.78 124.68 175.94 ;
      RECT 124.06 175.26 124.22 175.94 ;
      RECT 121.66 175.36 121.94 175.52 ;
      RECT 121.76 175.26 124.22 175.42 ;
      RECT 121.76 181.3 124.22 181.46 ;
      RECT 124.06 180.78 124.22 181.46 ;
      RECT 121.66 181.2 121.94 181.36 ;
      RECT 124.06 180.78 124.68 180.94 ;
      RECT 124.06 182.58 124.68 182.74 ;
      RECT 124.06 182.06 124.22 182.74 ;
      RECT 121.66 182.16 121.94 182.32 ;
      RECT 121.76 182.06 124.22 182.22 ;
      RECT 121.76 188.1 124.22 188.26 ;
      RECT 124.06 187.58 124.22 188.26 ;
      RECT 121.66 188 121.94 188.16 ;
      RECT 124.06 187.58 124.68 187.74 ;
      RECT 124.06 189.38 124.68 189.54 ;
      RECT 124.06 188.86 124.22 189.54 ;
      RECT 121.66 188.96 121.94 189.12 ;
      RECT 121.76 188.86 124.22 189.02 ;
      RECT 121.76 194.9 124.22 195.06 ;
      RECT 124.06 194.38 124.22 195.06 ;
      RECT 121.66 194.8 121.94 194.96 ;
      RECT 124.06 194.38 124.68 194.54 ;
      RECT 124.06 196.18 124.68 196.34 ;
      RECT 124.06 195.66 124.22 196.34 ;
      RECT 121.66 195.76 121.94 195.92 ;
      RECT 121.76 195.66 124.22 195.82 ;
      RECT 121.76 201.7 124.22 201.86 ;
      RECT 124.06 201.18 124.22 201.86 ;
      RECT 121.66 201.6 121.94 201.76 ;
      RECT 124.06 201.18 124.68 201.34 ;
      RECT 124.06 202.98 124.68 203.14 ;
      RECT 124.06 202.46 124.22 203.14 ;
      RECT 121.66 202.56 121.94 202.72 ;
      RECT 121.76 202.46 124.22 202.62 ;
      RECT 121.76 208.5 124.22 208.66 ;
      RECT 124.06 207.98 124.22 208.66 ;
      RECT 121.66 208.4 121.94 208.56 ;
      RECT 124.06 207.98 124.68 208.14 ;
      RECT 124.06 209.78 124.68 209.94 ;
      RECT 124.06 209.26 124.22 209.94 ;
      RECT 121.66 209.36 121.94 209.52 ;
      RECT 121.76 209.26 124.22 209.42 ;
      RECT 121.76 215.3 124.22 215.46 ;
      RECT 124.06 214.78 124.22 215.46 ;
      RECT 121.66 215.2 121.94 215.36 ;
      RECT 124.06 214.78 124.68 214.94 ;
      RECT 124.06 216.58 124.68 216.74 ;
      RECT 124.06 216.06 124.22 216.74 ;
      RECT 121.66 216.16 121.94 216.32 ;
      RECT 121.76 216.06 124.22 216.22 ;
      RECT 121.76 222.1 124.22 222.26 ;
      RECT 124.06 221.58 124.22 222.26 ;
      RECT 121.66 222 121.94 222.16 ;
      RECT 124.06 221.58 124.68 221.74 ;
      RECT 124.06 223.38 124.68 223.54 ;
      RECT 124.06 222.86 124.22 223.54 ;
      RECT 121.66 222.96 121.94 223.12 ;
      RECT 121.76 222.86 124.22 223.02 ;
      RECT 121.76 228.9 124.22 229.06 ;
      RECT 124.06 228.38 124.22 229.06 ;
      RECT 121.66 228.8 121.94 228.96 ;
      RECT 124.06 228.38 124.68 228.54 ;
      RECT 124.06 230.18 124.68 230.34 ;
      RECT 124.06 229.66 124.22 230.34 ;
      RECT 121.66 229.76 121.94 229.92 ;
      RECT 121.76 229.66 124.22 229.82 ;
      RECT 121.76 235.7 124.22 235.86 ;
      RECT 124.06 235.18 124.22 235.86 ;
      RECT 121.66 235.6 121.94 235.76 ;
      RECT 124.06 235.18 124.68 235.34 ;
      RECT 124.06 236.98 124.68 237.14 ;
      RECT 124.06 236.46 124.22 237.14 ;
      RECT 121.66 236.56 121.94 236.72 ;
      RECT 121.76 236.46 124.22 236.62 ;
      RECT 121.76 242.5 124.22 242.66 ;
      RECT 124.06 241.98 124.22 242.66 ;
      RECT 121.66 242.4 121.94 242.56 ;
      RECT 124.06 241.98 124.68 242.14 ;
      RECT 124.06 243.78 124.68 243.94 ;
      RECT 124.06 243.26 124.22 243.94 ;
      RECT 121.66 243.36 121.94 243.52 ;
      RECT 121.76 243.26 124.22 243.42 ;
      RECT 121.76 249.3 124.22 249.46 ;
      RECT 124.06 248.78 124.22 249.46 ;
      RECT 121.66 249.2 121.94 249.36 ;
      RECT 124.06 248.78 124.68 248.94 ;
      RECT 124.06 250.58 124.68 250.74 ;
      RECT 124.06 250.06 124.22 250.74 ;
      RECT 121.66 250.16 121.94 250.32 ;
      RECT 121.76 250.06 124.22 250.22 ;
      RECT 121.76 256.1 124.22 256.26 ;
      RECT 124.06 255.58 124.22 256.26 ;
      RECT 121.66 256 121.94 256.16 ;
      RECT 124.06 255.58 124.68 255.74 ;
      RECT 124.06 257.38 124.68 257.54 ;
      RECT 124.06 256.86 124.22 257.54 ;
      RECT 121.66 256.96 121.94 257.12 ;
      RECT 121.76 256.86 124.22 257.02 ;
      RECT 121.76 262.9 124.22 263.06 ;
      RECT 124.06 262.38 124.22 263.06 ;
      RECT 121.66 262.8 121.94 262.96 ;
      RECT 124.06 262.38 124.68 262.54 ;
      RECT 124.06 264.18 124.68 264.34 ;
      RECT 124.06 263.66 124.22 264.34 ;
      RECT 121.66 263.76 121.94 263.92 ;
      RECT 121.76 263.66 124.22 263.82 ;
      RECT 121.76 269.7 124.22 269.86 ;
      RECT 124.06 269.18 124.22 269.86 ;
      RECT 121.66 269.6 121.94 269.76 ;
      RECT 124.06 269.18 124.68 269.34 ;
      RECT 124.06 270.98 124.68 271.14 ;
      RECT 124.06 270.46 124.22 271.14 ;
      RECT 121.66 270.56 121.94 270.72 ;
      RECT 121.76 270.46 124.22 270.62 ;
      RECT 121.76 276.5 124.22 276.66 ;
      RECT 124.06 275.98 124.22 276.66 ;
      RECT 121.66 276.4 121.94 276.56 ;
      RECT 124.06 275.98 124.68 276.14 ;
      RECT 124.06 277.78 124.68 277.94 ;
      RECT 124.06 277.26 124.22 277.94 ;
      RECT 121.66 277.36 121.94 277.52 ;
      RECT 121.76 277.26 124.22 277.42 ;
      RECT 121.76 283.3 124.22 283.46 ;
      RECT 124.06 282.78 124.22 283.46 ;
      RECT 121.66 283.2 121.94 283.36 ;
      RECT 124.06 282.78 124.68 282.94 ;
      RECT 124.06 284.58 124.68 284.74 ;
      RECT 124.06 284.06 124.22 284.74 ;
      RECT 121.66 284.16 121.94 284.32 ;
      RECT 121.76 284.06 124.22 284.22 ;
      RECT 121.76 290.1 124.22 290.26 ;
      RECT 124.06 289.58 124.22 290.26 ;
      RECT 121.66 290 121.94 290.16 ;
      RECT 124.06 289.58 124.68 289.74 ;
      RECT 124.06 291.38 124.68 291.54 ;
      RECT 124.06 290.86 124.22 291.54 ;
      RECT 121.66 290.96 121.94 291.12 ;
      RECT 121.76 290.86 124.22 291.02 ;
      RECT 121.76 296.9 124.22 297.06 ;
      RECT 124.06 296.38 124.22 297.06 ;
      RECT 121.66 296.8 121.94 296.96 ;
      RECT 124.06 296.38 124.68 296.54 ;
      RECT 124.06 298.18 124.68 298.34 ;
      RECT 124.06 297.66 124.22 298.34 ;
      RECT 121.66 297.76 121.94 297.92 ;
      RECT 121.76 297.66 124.22 297.82 ;
      RECT 121.76 303.7 124.22 303.86 ;
      RECT 124.06 303.18 124.22 303.86 ;
      RECT 121.66 303.6 121.94 303.76 ;
      RECT 124.06 303.18 124.68 303.34 ;
      RECT 124.06 304.98 124.68 305.14 ;
      RECT 124.06 304.46 124.22 305.14 ;
      RECT 121.66 304.56 121.94 304.72 ;
      RECT 121.76 304.46 124.22 304.62 ;
      RECT 121.76 310.5 124.22 310.66 ;
      RECT 124.06 309.98 124.22 310.66 ;
      RECT 121.66 310.4 121.94 310.56 ;
      RECT 124.06 309.98 124.68 310.14 ;
      RECT 124.06 311.78 124.68 311.94 ;
      RECT 124.06 311.26 124.22 311.94 ;
      RECT 121.66 311.36 121.94 311.52 ;
      RECT 121.76 311.26 124.22 311.42 ;
      RECT 121.76 317.3 124.22 317.46 ;
      RECT 124.06 316.78 124.22 317.46 ;
      RECT 121.66 317.2 121.94 317.36 ;
      RECT 124.06 316.78 124.68 316.94 ;
      RECT 124.06 318.58 124.68 318.74 ;
      RECT 124.06 318.06 124.22 318.74 ;
      RECT 121.66 318.16 121.94 318.32 ;
      RECT 121.76 318.06 124.22 318.22 ;
      RECT 121.76 324.1 124.22 324.26 ;
      RECT 124.06 323.58 124.22 324.26 ;
      RECT 121.66 324 121.94 324.16 ;
      RECT 124.06 323.58 124.68 323.74 ;
      RECT 124.06 325.38 124.68 325.54 ;
      RECT 124.06 324.86 124.22 325.54 ;
      RECT 121.66 324.96 121.94 325.12 ;
      RECT 121.76 324.86 124.22 325.02 ;
      RECT 121.76 330.9 124.22 331.06 ;
      RECT 124.06 330.38 124.22 331.06 ;
      RECT 121.66 330.8 121.94 330.96 ;
      RECT 124.06 330.38 124.68 330.54 ;
      RECT 124.06 332.18 124.68 332.34 ;
      RECT 124.06 331.66 124.22 332.34 ;
      RECT 121.66 331.76 121.94 331.92 ;
      RECT 121.76 331.66 124.22 331.82 ;
      RECT 121.76 337.7 124.22 337.86 ;
      RECT 124.06 337.18 124.22 337.86 ;
      RECT 121.66 337.6 121.94 337.76 ;
      RECT 124.06 337.18 124.68 337.34 ;
      RECT 124.06 338.98 124.68 339.14 ;
      RECT 124.06 338.46 124.22 339.14 ;
      RECT 121.66 338.56 121.94 338.72 ;
      RECT 121.76 338.46 124.22 338.62 ;
      RECT 121.76 344.5 124.22 344.66 ;
      RECT 124.06 343.98 124.22 344.66 ;
      RECT 121.66 344.4 121.94 344.56 ;
      RECT 124.06 343.98 124.68 344.14 ;
      RECT 124.06 345.78 124.68 345.94 ;
      RECT 124.06 345.26 124.22 345.94 ;
      RECT 121.66 345.36 121.94 345.52 ;
      RECT 121.76 345.26 124.22 345.42 ;
      RECT 121.76 351.3 124.22 351.46 ;
      RECT 124.06 350.78 124.22 351.46 ;
      RECT 121.66 351.2 121.94 351.36 ;
      RECT 124.06 350.78 124.68 350.94 ;
      RECT 124.06 352.58 124.68 352.74 ;
      RECT 124.06 352.06 124.22 352.74 ;
      RECT 121.66 352.16 121.94 352.32 ;
      RECT 121.76 352.06 124.22 352.22 ;
      RECT 121.76 358.1 124.22 358.26 ;
      RECT 124.06 357.58 124.22 358.26 ;
      RECT 121.66 358 121.94 358.16 ;
      RECT 124.06 357.58 124.68 357.74 ;
      RECT 124.06 359.38 124.68 359.54 ;
      RECT 124.06 358.86 124.22 359.54 ;
      RECT 121.66 358.96 121.94 359.12 ;
      RECT 121.76 358.86 124.22 359.02 ;
      RECT 121.76 364.9 124.22 365.06 ;
      RECT 124.06 364.38 124.22 365.06 ;
      RECT 121.66 364.8 121.94 364.96 ;
      RECT 124.06 364.38 124.68 364.54 ;
      RECT 124.06 366.18 124.68 366.34 ;
      RECT 124.06 365.66 124.22 366.34 ;
      RECT 121.66 365.76 121.94 365.92 ;
      RECT 121.76 365.66 124.22 365.82 ;
      RECT 121.76 371.7 124.22 371.86 ;
      RECT 124.06 371.18 124.22 371.86 ;
      RECT 121.66 371.6 121.94 371.76 ;
      RECT 124.06 371.18 124.68 371.34 ;
      RECT 124.06 372.98 124.68 373.14 ;
      RECT 124.06 372.46 124.22 373.14 ;
      RECT 121.66 372.56 121.94 372.72 ;
      RECT 121.76 372.46 124.22 372.62 ;
      RECT 121.76 378.5 124.22 378.66 ;
      RECT 124.06 377.98 124.22 378.66 ;
      RECT 121.66 378.4 121.94 378.56 ;
      RECT 124.06 377.98 124.68 378.14 ;
      RECT 124.06 379.78 124.68 379.94 ;
      RECT 124.06 379.26 124.22 379.94 ;
      RECT 121.66 379.36 121.94 379.52 ;
      RECT 121.76 379.26 124.22 379.42 ;
      RECT 121.76 385.3 124.22 385.46 ;
      RECT 124.06 384.78 124.22 385.46 ;
      RECT 121.66 385.2 121.94 385.36 ;
      RECT 124.06 384.78 124.68 384.94 ;
      RECT 124.06 386.58 124.68 386.74 ;
      RECT 124.06 386.06 124.22 386.74 ;
      RECT 121.66 386.16 121.94 386.32 ;
      RECT 121.76 386.06 124.22 386.22 ;
      RECT 121.76 392.1 124.22 392.26 ;
      RECT 124.06 391.58 124.22 392.26 ;
      RECT 121.66 392 121.94 392.16 ;
      RECT 124.06 391.58 124.68 391.74 ;
      RECT 124.06 393.38 124.68 393.54 ;
      RECT 124.06 392.86 124.22 393.54 ;
      RECT 121.66 392.96 121.94 393.12 ;
      RECT 121.76 392.86 124.22 393.02 ;
      RECT 121.76 398.9 124.22 399.06 ;
      RECT 124.06 398.38 124.22 399.06 ;
      RECT 121.66 398.8 121.94 398.96 ;
      RECT 124.06 398.38 124.68 398.54 ;
      RECT 124.06 400.18 124.68 400.34 ;
      RECT 124.06 399.66 124.22 400.34 ;
      RECT 121.66 399.76 121.94 399.92 ;
      RECT 121.76 399.66 124.22 399.82 ;
      RECT 121.76 405.7 124.22 405.86 ;
      RECT 124.06 405.18 124.22 405.86 ;
      RECT 121.66 405.6 121.94 405.76 ;
      RECT 124.06 405.18 124.68 405.34 ;
      RECT 124.06 406.98 124.68 407.14 ;
      RECT 124.06 406.46 124.22 407.14 ;
      RECT 121.66 406.56 121.94 406.72 ;
      RECT 121.76 406.46 124.22 406.62 ;
      RECT 121.76 412.5 124.22 412.66 ;
      RECT 124.06 411.98 124.22 412.66 ;
      RECT 121.66 412.4 121.94 412.56 ;
      RECT 124.06 411.98 124.68 412.14 ;
      RECT 124.06 413.78 124.68 413.94 ;
      RECT 124.06 413.26 124.22 413.94 ;
      RECT 121.66 413.36 121.94 413.52 ;
      RECT 121.76 413.26 124.22 413.42 ;
      RECT 121.76 419.3 124.22 419.46 ;
      RECT 124.06 418.78 124.22 419.46 ;
      RECT 121.66 419.2 121.94 419.36 ;
      RECT 124.06 418.78 124.68 418.94 ;
      RECT 124.06 420.58 124.68 420.74 ;
      RECT 124.06 420.06 124.22 420.74 ;
      RECT 121.66 420.16 121.94 420.32 ;
      RECT 121.76 420.06 124.22 420.22 ;
      RECT 121.76 426.1 124.22 426.26 ;
      RECT 124.06 425.58 124.22 426.26 ;
      RECT 121.66 426 121.94 426.16 ;
      RECT 124.06 425.58 124.68 425.74 ;
      RECT 124.06 427.38 124.68 427.54 ;
      RECT 124.06 426.86 124.22 427.54 ;
      RECT 121.66 426.96 121.94 427.12 ;
      RECT 121.76 426.86 124.22 427.02 ;
      RECT 121.76 432.9 124.22 433.06 ;
      RECT 124.06 432.38 124.22 433.06 ;
      RECT 121.66 432.8 121.94 432.96 ;
      RECT 124.06 432.38 124.68 432.54 ;
      RECT 124.06 434.18 124.68 434.34 ;
      RECT 124.06 433.66 124.22 434.34 ;
      RECT 121.66 433.76 121.94 433.92 ;
      RECT 121.76 433.66 124.22 433.82 ;
      RECT 121.76 439.7 124.22 439.86 ;
      RECT 124.06 439.18 124.22 439.86 ;
      RECT 121.66 439.6 121.94 439.76 ;
      RECT 124.06 439.18 124.68 439.34 ;
      RECT 124.06 440.98 124.68 441.14 ;
      RECT 124.06 440.46 124.22 441.14 ;
      RECT 121.66 440.56 121.94 440.72 ;
      RECT 121.76 440.46 124.22 440.62 ;
      RECT 121.76 446.5 124.22 446.66 ;
      RECT 124.06 445.98 124.22 446.66 ;
      RECT 121.66 446.4 121.94 446.56 ;
      RECT 124.06 445.98 124.68 446.14 ;
      RECT 124.06 447.78 124.68 447.94 ;
      RECT 124.06 447.26 124.22 447.94 ;
      RECT 121.66 447.36 121.94 447.52 ;
      RECT 121.76 447.26 124.22 447.42 ;
      RECT 121.76 453.3 124.22 453.46 ;
      RECT 124.06 452.78 124.22 453.46 ;
      RECT 121.66 453.2 121.94 453.36 ;
      RECT 124.06 452.78 124.68 452.94 ;
      RECT 124.06 454.58 124.68 454.74 ;
      RECT 124.06 454.06 124.22 454.74 ;
      RECT 121.66 454.16 121.94 454.32 ;
      RECT 121.76 454.06 124.22 454.22 ;
      RECT 121.76 460.1 124.22 460.26 ;
      RECT 124.06 459.58 124.22 460.26 ;
      RECT 121.66 460 121.94 460.16 ;
      RECT 124.06 459.58 124.68 459.74 ;
      RECT 124.06 461.38 124.68 461.54 ;
      RECT 124.06 460.86 124.22 461.54 ;
      RECT 121.66 460.96 121.94 461.12 ;
      RECT 121.76 460.86 124.22 461.02 ;
      RECT 121.76 466.9 124.22 467.06 ;
      RECT 124.06 466.38 124.22 467.06 ;
      RECT 121.66 466.8 121.94 466.96 ;
      RECT 124.06 466.38 124.68 466.54 ;
      RECT 124.06 468.18 124.68 468.34 ;
      RECT 124.06 467.66 124.22 468.34 ;
      RECT 121.66 467.76 121.94 467.92 ;
      RECT 121.76 467.66 124.22 467.82 ;
      RECT 121.76 473.7 124.22 473.86 ;
      RECT 124.06 473.18 124.22 473.86 ;
      RECT 121.66 473.6 121.94 473.76 ;
      RECT 124.06 473.18 124.68 473.34 ;
      RECT 124.06 474.98 124.68 475.14 ;
      RECT 124.06 474.46 124.22 475.14 ;
      RECT 121.66 474.56 121.94 474.72 ;
      RECT 121.76 474.46 124.22 474.62 ;
      RECT 121.76 480.5 124.22 480.66 ;
      RECT 124.06 479.98 124.22 480.66 ;
      RECT 121.66 480.4 121.94 480.56 ;
      RECT 124.06 479.98 124.68 480.14 ;
      RECT 124.06 481.78 124.68 481.94 ;
      RECT 124.06 481.26 124.22 481.94 ;
      RECT 121.66 481.36 121.94 481.52 ;
      RECT 121.76 481.26 124.22 481.42 ;
      RECT 121.76 487.3 124.22 487.46 ;
      RECT 124.06 486.78 124.22 487.46 ;
      RECT 121.66 487.2 121.94 487.36 ;
      RECT 124.06 486.78 124.68 486.94 ;
      RECT 124.06 488.58 124.68 488.74 ;
      RECT 124.06 488.06 124.22 488.74 ;
      RECT 121.66 488.16 121.94 488.32 ;
      RECT 121.76 488.06 124.22 488.22 ;
      RECT 121.76 494.1 124.22 494.26 ;
      RECT 124.06 493.58 124.22 494.26 ;
      RECT 121.66 494 121.94 494.16 ;
      RECT 124.06 493.58 124.68 493.74 ;
      RECT 124.06 495.38 124.68 495.54 ;
      RECT 124.06 494.86 124.22 495.54 ;
      RECT 121.66 494.96 121.94 495.12 ;
      RECT 121.76 494.86 124.22 495.02 ;
      RECT 121.76 500.9 124.22 501.06 ;
      RECT 124.06 500.38 124.22 501.06 ;
      RECT 121.66 500.8 121.94 500.96 ;
      RECT 124.06 500.38 124.68 500.54 ;
      RECT 124.06 502.18 124.68 502.34 ;
      RECT 124.06 501.66 124.22 502.34 ;
      RECT 121.66 501.76 121.94 501.92 ;
      RECT 121.76 501.66 124.22 501.82 ;
      RECT 121.62 506.12 121.78 507.58 ;
      RECT 121.62 506.12 124.62 506.28 ;
      RECT 123.95 31.09 124.11 35.75 ;
      RECT 123.85 32.25 124.11 32.53 ;
      RECT 123.91 49.75 124.11 51.3 ;
      RECT 123.95 46.54 124.11 51.3 ;
      RECT 123.51 49.6 123.67 51.7 ;
      RECT 123.07 49.6 123.67 49.76 ;
      RECT 123.07 32.06 123.23 49.76 ;
      RECT 123.07 45.9 123.89 46.06 ;
      RECT 123.07 36.23 123.89 36.39 ;
      RECT 123.07 32.06 123.67 32.22 ;
      RECT 123.51 30.54 123.67 32.22 ;
      RECT 123.18 70.38 123.88 70.54 ;
      RECT 123.24 70.18 123.6 70.54 ;
      RECT 123.24 71.98 123.6 72.34 ;
      RECT 123.18 71.98 123.88 72.14 ;
      RECT 123.18 73.78 123.88 73.94 ;
      RECT 123.24 73.58 123.6 73.94 ;
      RECT 123.24 75.38 123.6 75.74 ;
      RECT 123.18 75.38 123.88 75.54 ;
      RECT 123.18 77.18 123.88 77.34 ;
      RECT 123.24 76.98 123.6 77.34 ;
      RECT 123.24 78.78 123.6 79.14 ;
      RECT 123.18 78.78 123.88 78.94 ;
      RECT 123.18 80.58 123.88 80.74 ;
      RECT 123.24 80.38 123.6 80.74 ;
      RECT 123.24 82.18 123.6 82.54 ;
      RECT 123.18 82.18 123.88 82.34 ;
      RECT 123.18 83.98 123.88 84.14 ;
      RECT 123.24 83.78 123.6 84.14 ;
      RECT 123.24 85.58 123.6 85.94 ;
      RECT 123.18 85.58 123.88 85.74 ;
      RECT 123.18 87.38 123.88 87.54 ;
      RECT 123.24 87.18 123.6 87.54 ;
      RECT 123.24 88.98 123.6 89.34 ;
      RECT 123.18 88.98 123.88 89.14 ;
      RECT 123.18 90.78 123.88 90.94 ;
      RECT 123.24 90.58 123.6 90.94 ;
      RECT 123.24 92.38 123.6 92.74 ;
      RECT 123.18 92.38 123.88 92.54 ;
      RECT 123.18 94.18 123.88 94.34 ;
      RECT 123.24 93.98 123.6 94.34 ;
      RECT 123.24 95.78 123.6 96.14 ;
      RECT 123.18 95.78 123.88 95.94 ;
      RECT 123.18 97.58 123.88 97.74 ;
      RECT 123.24 97.38 123.6 97.74 ;
      RECT 123.24 99.18 123.6 99.54 ;
      RECT 123.18 99.18 123.88 99.34 ;
      RECT 123.18 100.98 123.88 101.14 ;
      RECT 123.24 100.78 123.6 101.14 ;
      RECT 123.24 102.58 123.6 102.94 ;
      RECT 123.18 102.58 123.88 102.74 ;
      RECT 123.18 104.38 123.88 104.54 ;
      RECT 123.24 104.18 123.6 104.54 ;
      RECT 123.24 105.98 123.6 106.34 ;
      RECT 123.18 105.98 123.88 106.14 ;
      RECT 123.18 107.78 123.88 107.94 ;
      RECT 123.24 107.58 123.6 107.94 ;
      RECT 123.24 109.38 123.6 109.74 ;
      RECT 123.18 109.38 123.88 109.54 ;
      RECT 123.18 111.18 123.88 111.34 ;
      RECT 123.24 110.98 123.6 111.34 ;
      RECT 123.24 112.78 123.6 113.14 ;
      RECT 123.18 112.78 123.88 112.94 ;
      RECT 123.18 114.58 123.88 114.74 ;
      RECT 123.24 114.38 123.6 114.74 ;
      RECT 123.24 116.18 123.6 116.54 ;
      RECT 123.18 116.18 123.88 116.34 ;
      RECT 123.18 117.98 123.88 118.14 ;
      RECT 123.24 117.78 123.6 118.14 ;
      RECT 123.24 119.58 123.6 119.94 ;
      RECT 123.18 119.58 123.88 119.74 ;
      RECT 123.18 121.38 123.88 121.54 ;
      RECT 123.24 121.18 123.6 121.54 ;
      RECT 123.24 122.98 123.6 123.34 ;
      RECT 123.18 122.98 123.88 123.14 ;
      RECT 123.18 124.78 123.88 124.94 ;
      RECT 123.24 124.58 123.6 124.94 ;
      RECT 123.24 126.38 123.6 126.74 ;
      RECT 123.18 126.38 123.88 126.54 ;
      RECT 123.18 128.18 123.88 128.34 ;
      RECT 123.24 127.98 123.6 128.34 ;
      RECT 123.24 129.78 123.6 130.14 ;
      RECT 123.18 129.78 123.88 129.94 ;
      RECT 123.18 131.58 123.88 131.74 ;
      RECT 123.24 131.38 123.6 131.74 ;
      RECT 123.24 133.18 123.6 133.54 ;
      RECT 123.18 133.18 123.88 133.34 ;
      RECT 123.18 134.98 123.88 135.14 ;
      RECT 123.24 134.78 123.6 135.14 ;
      RECT 123.24 136.58 123.6 136.94 ;
      RECT 123.18 136.58 123.88 136.74 ;
      RECT 123.18 138.38 123.88 138.54 ;
      RECT 123.24 138.18 123.6 138.54 ;
      RECT 123.24 139.98 123.6 140.34 ;
      RECT 123.18 139.98 123.88 140.14 ;
      RECT 123.18 141.78 123.88 141.94 ;
      RECT 123.24 141.58 123.6 141.94 ;
      RECT 123.24 143.38 123.6 143.74 ;
      RECT 123.18 143.38 123.88 143.54 ;
      RECT 123.18 145.18 123.88 145.34 ;
      RECT 123.24 144.98 123.6 145.34 ;
      RECT 123.24 146.78 123.6 147.14 ;
      RECT 123.18 146.78 123.88 146.94 ;
      RECT 123.18 148.58 123.88 148.74 ;
      RECT 123.24 148.38 123.6 148.74 ;
      RECT 123.24 150.18 123.6 150.54 ;
      RECT 123.18 150.18 123.88 150.34 ;
      RECT 123.18 151.98 123.88 152.14 ;
      RECT 123.24 151.78 123.6 152.14 ;
      RECT 123.24 153.58 123.6 153.94 ;
      RECT 123.18 153.58 123.88 153.74 ;
      RECT 123.18 155.38 123.88 155.54 ;
      RECT 123.24 155.18 123.6 155.54 ;
      RECT 123.24 156.98 123.6 157.34 ;
      RECT 123.18 156.98 123.88 157.14 ;
      RECT 123.18 158.78 123.88 158.94 ;
      RECT 123.24 158.58 123.6 158.94 ;
      RECT 123.24 160.38 123.6 160.74 ;
      RECT 123.18 160.38 123.88 160.54 ;
      RECT 123.18 162.18 123.88 162.34 ;
      RECT 123.24 161.98 123.6 162.34 ;
      RECT 123.24 163.78 123.6 164.14 ;
      RECT 123.18 163.78 123.88 163.94 ;
      RECT 123.18 165.58 123.88 165.74 ;
      RECT 123.24 165.38 123.6 165.74 ;
      RECT 123.24 167.18 123.6 167.54 ;
      RECT 123.18 167.18 123.88 167.34 ;
      RECT 123.18 168.98 123.88 169.14 ;
      RECT 123.24 168.78 123.6 169.14 ;
      RECT 123.24 170.58 123.6 170.94 ;
      RECT 123.18 170.58 123.88 170.74 ;
      RECT 123.18 172.38 123.88 172.54 ;
      RECT 123.24 172.18 123.6 172.54 ;
      RECT 123.24 173.98 123.6 174.34 ;
      RECT 123.18 173.98 123.88 174.14 ;
      RECT 123.18 175.78 123.88 175.94 ;
      RECT 123.24 175.58 123.6 175.94 ;
      RECT 123.24 177.38 123.6 177.74 ;
      RECT 123.18 177.38 123.88 177.54 ;
      RECT 123.18 179.18 123.88 179.34 ;
      RECT 123.24 178.98 123.6 179.34 ;
      RECT 123.24 180.78 123.6 181.14 ;
      RECT 123.18 180.78 123.88 180.94 ;
      RECT 123.18 182.58 123.88 182.74 ;
      RECT 123.24 182.38 123.6 182.74 ;
      RECT 123.24 184.18 123.6 184.54 ;
      RECT 123.18 184.18 123.88 184.34 ;
      RECT 123.18 185.98 123.88 186.14 ;
      RECT 123.24 185.78 123.6 186.14 ;
      RECT 123.24 187.58 123.6 187.94 ;
      RECT 123.18 187.58 123.88 187.74 ;
      RECT 123.18 189.38 123.88 189.54 ;
      RECT 123.24 189.18 123.6 189.54 ;
      RECT 123.24 190.98 123.6 191.34 ;
      RECT 123.18 190.98 123.88 191.14 ;
      RECT 123.18 192.78 123.88 192.94 ;
      RECT 123.24 192.58 123.6 192.94 ;
      RECT 123.24 194.38 123.6 194.74 ;
      RECT 123.18 194.38 123.88 194.54 ;
      RECT 123.18 196.18 123.88 196.34 ;
      RECT 123.24 195.98 123.6 196.34 ;
      RECT 123.24 197.78 123.6 198.14 ;
      RECT 123.18 197.78 123.88 197.94 ;
      RECT 123.18 199.58 123.88 199.74 ;
      RECT 123.24 199.38 123.6 199.74 ;
      RECT 123.24 201.18 123.6 201.54 ;
      RECT 123.18 201.18 123.88 201.34 ;
      RECT 123.18 202.98 123.88 203.14 ;
      RECT 123.24 202.78 123.6 203.14 ;
      RECT 123.24 204.58 123.6 204.94 ;
      RECT 123.18 204.58 123.88 204.74 ;
      RECT 123.18 206.38 123.88 206.54 ;
      RECT 123.24 206.18 123.6 206.54 ;
      RECT 123.24 207.98 123.6 208.34 ;
      RECT 123.18 207.98 123.88 208.14 ;
      RECT 123.18 209.78 123.88 209.94 ;
      RECT 123.24 209.58 123.6 209.94 ;
      RECT 123.24 211.38 123.6 211.74 ;
      RECT 123.18 211.38 123.88 211.54 ;
      RECT 123.18 213.18 123.88 213.34 ;
      RECT 123.24 212.98 123.6 213.34 ;
      RECT 123.24 214.78 123.6 215.14 ;
      RECT 123.18 214.78 123.88 214.94 ;
      RECT 123.18 216.58 123.88 216.74 ;
      RECT 123.24 216.38 123.6 216.74 ;
      RECT 123.24 218.18 123.6 218.54 ;
      RECT 123.18 218.18 123.88 218.34 ;
      RECT 123.18 219.98 123.88 220.14 ;
      RECT 123.24 219.78 123.6 220.14 ;
      RECT 123.24 221.58 123.6 221.94 ;
      RECT 123.18 221.58 123.88 221.74 ;
      RECT 123.18 223.38 123.88 223.54 ;
      RECT 123.24 223.18 123.6 223.54 ;
      RECT 123.24 224.98 123.6 225.34 ;
      RECT 123.18 224.98 123.88 225.14 ;
      RECT 123.18 226.78 123.88 226.94 ;
      RECT 123.24 226.58 123.6 226.94 ;
      RECT 123.24 228.38 123.6 228.74 ;
      RECT 123.18 228.38 123.88 228.54 ;
      RECT 123.18 230.18 123.88 230.34 ;
      RECT 123.24 229.98 123.6 230.34 ;
      RECT 123.24 231.78 123.6 232.14 ;
      RECT 123.18 231.78 123.88 231.94 ;
      RECT 123.18 233.58 123.88 233.74 ;
      RECT 123.24 233.38 123.6 233.74 ;
      RECT 123.24 235.18 123.6 235.54 ;
      RECT 123.18 235.18 123.88 235.34 ;
      RECT 123.18 236.98 123.88 237.14 ;
      RECT 123.24 236.78 123.6 237.14 ;
      RECT 123.24 238.58 123.6 238.94 ;
      RECT 123.18 238.58 123.88 238.74 ;
      RECT 123.18 240.38 123.88 240.54 ;
      RECT 123.24 240.18 123.6 240.54 ;
      RECT 123.24 241.98 123.6 242.34 ;
      RECT 123.18 241.98 123.88 242.14 ;
      RECT 123.18 243.78 123.88 243.94 ;
      RECT 123.24 243.58 123.6 243.94 ;
      RECT 123.24 245.38 123.6 245.74 ;
      RECT 123.18 245.38 123.88 245.54 ;
      RECT 123.18 247.18 123.88 247.34 ;
      RECT 123.24 246.98 123.6 247.34 ;
      RECT 123.24 248.78 123.6 249.14 ;
      RECT 123.18 248.78 123.88 248.94 ;
      RECT 123.18 250.58 123.88 250.74 ;
      RECT 123.24 250.38 123.6 250.74 ;
      RECT 123.24 252.18 123.6 252.54 ;
      RECT 123.18 252.18 123.88 252.34 ;
      RECT 123.18 253.98 123.88 254.14 ;
      RECT 123.24 253.78 123.6 254.14 ;
      RECT 123.24 255.58 123.6 255.94 ;
      RECT 123.18 255.58 123.88 255.74 ;
      RECT 123.18 257.38 123.88 257.54 ;
      RECT 123.24 257.18 123.6 257.54 ;
      RECT 123.24 258.98 123.6 259.34 ;
      RECT 123.18 258.98 123.88 259.14 ;
      RECT 123.18 260.78 123.88 260.94 ;
      RECT 123.24 260.58 123.6 260.94 ;
      RECT 123.24 262.38 123.6 262.74 ;
      RECT 123.18 262.38 123.88 262.54 ;
      RECT 123.18 264.18 123.88 264.34 ;
      RECT 123.24 263.98 123.6 264.34 ;
      RECT 123.24 265.78 123.6 266.14 ;
      RECT 123.18 265.78 123.88 265.94 ;
      RECT 123.18 267.58 123.88 267.74 ;
      RECT 123.24 267.38 123.6 267.74 ;
      RECT 123.24 269.18 123.6 269.54 ;
      RECT 123.18 269.18 123.88 269.34 ;
      RECT 123.18 270.98 123.88 271.14 ;
      RECT 123.24 270.78 123.6 271.14 ;
      RECT 123.24 272.58 123.6 272.94 ;
      RECT 123.18 272.58 123.88 272.74 ;
      RECT 123.18 274.38 123.88 274.54 ;
      RECT 123.24 274.18 123.6 274.54 ;
      RECT 123.24 275.98 123.6 276.34 ;
      RECT 123.18 275.98 123.88 276.14 ;
      RECT 123.18 277.78 123.88 277.94 ;
      RECT 123.24 277.58 123.6 277.94 ;
      RECT 123.24 279.38 123.6 279.74 ;
      RECT 123.18 279.38 123.88 279.54 ;
      RECT 123.18 281.18 123.88 281.34 ;
      RECT 123.24 280.98 123.6 281.34 ;
      RECT 123.24 282.78 123.6 283.14 ;
      RECT 123.18 282.78 123.88 282.94 ;
      RECT 123.18 284.58 123.88 284.74 ;
      RECT 123.24 284.38 123.6 284.74 ;
      RECT 123.24 286.18 123.6 286.54 ;
      RECT 123.18 286.18 123.88 286.34 ;
      RECT 123.18 287.98 123.88 288.14 ;
      RECT 123.24 287.78 123.6 288.14 ;
      RECT 123.24 289.58 123.6 289.94 ;
      RECT 123.18 289.58 123.88 289.74 ;
      RECT 123.18 291.38 123.88 291.54 ;
      RECT 123.24 291.18 123.6 291.54 ;
      RECT 123.24 292.98 123.6 293.34 ;
      RECT 123.18 292.98 123.88 293.14 ;
      RECT 123.18 294.78 123.88 294.94 ;
      RECT 123.24 294.58 123.6 294.94 ;
      RECT 123.24 296.38 123.6 296.74 ;
      RECT 123.18 296.38 123.88 296.54 ;
      RECT 123.18 298.18 123.88 298.34 ;
      RECT 123.24 297.98 123.6 298.34 ;
      RECT 123.24 299.78 123.6 300.14 ;
      RECT 123.18 299.78 123.88 299.94 ;
      RECT 123.18 301.58 123.88 301.74 ;
      RECT 123.24 301.38 123.6 301.74 ;
      RECT 123.24 303.18 123.6 303.54 ;
      RECT 123.18 303.18 123.88 303.34 ;
      RECT 123.18 304.98 123.88 305.14 ;
      RECT 123.24 304.78 123.6 305.14 ;
      RECT 123.24 306.58 123.6 306.94 ;
      RECT 123.18 306.58 123.88 306.74 ;
      RECT 123.18 308.38 123.88 308.54 ;
      RECT 123.24 308.18 123.6 308.54 ;
      RECT 123.24 309.98 123.6 310.34 ;
      RECT 123.18 309.98 123.88 310.14 ;
      RECT 123.18 311.78 123.88 311.94 ;
      RECT 123.24 311.58 123.6 311.94 ;
      RECT 123.24 313.38 123.6 313.74 ;
      RECT 123.18 313.38 123.88 313.54 ;
      RECT 123.18 315.18 123.88 315.34 ;
      RECT 123.24 314.98 123.6 315.34 ;
      RECT 123.24 316.78 123.6 317.14 ;
      RECT 123.18 316.78 123.88 316.94 ;
      RECT 123.18 318.58 123.88 318.74 ;
      RECT 123.24 318.38 123.6 318.74 ;
      RECT 123.24 320.18 123.6 320.54 ;
      RECT 123.18 320.18 123.88 320.34 ;
      RECT 123.18 321.98 123.88 322.14 ;
      RECT 123.24 321.78 123.6 322.14 ;
      RECT 123.24 323.58 123.6 323.94 ;
      RECT 123.18 323.58 123.88 323.74 ;
      RECT 123.18 325.38 123.88 325.54 ;
      RECT 123.24 325.18 123.6 325.54 ;
      RECT 123.24 326.98 123.6 327.34 ;
      RECT 123.18 326.98 123.88 327.14 ;
      RECT 123.18 328.78 123.88 328.94 ;
      RECT 123.24 328.58 123.6 328.94 ;
      RECT 123.24 330.38 123.6 330.74 ;
      RECT 123.18 330.38 123.88 330.54 ;
      RECT 123.18 332.18 123.88 332.34 ;
      RECT 123.24 331.98 123.6 332.34 ;
      RECT 123.24 333.78 123.6 334.14 ;
      RECT 123.18 333.78 123.88 333.94 ;
      RECT 123.18 335.58 123.88 335.74 ;
      RECT 123.24 335.38 123.6 335.74 ;
      RECT 123.24 337.18 123.6 337.54 ;
      RECT 123.18 337.18 123.88 337.34 ;
      RECT 123.18 338.98 123.88 339.14 ;
      RECT 123.24 338.78 123.6 339.14 ;
      RECT 123.24 340.58 123.6 340.94 ;
      RECT 123.18 340.58 123.88 340.74 ;
      RECT 123.18 342.38 123.88 342.54 ;
      RECT 123.24 342.18 123.6 342.54 ;
      RECT 123.24 343.98 123.6 344.34 ;
      RECT 123.18 343.98 123.88 344.14 ;
      RECT 123.18 345.78 123.88 345.94 ;
      RECT 123.24 345.58 123.6 345.94 ;
      RECT 123.24 347.38 123.6 347.74 ;
      RECT 123.18 347.38 123.88 347.54 ;
      RECT 123.18 349.18 123.88 349.34 ;
      RECT 123.24 348.98 123.6 349.34 ;
      RECT 123.24 350.78 123.6 351.14 ;
      RECT 123.18 350.78 123.88 350.94 ;
      RECT 123.18 352.58 123.88 352.74 ;
      RECT 123.24 352.38 123.6 352.74 ;
      RECT 123.24 354.18 123.6 354.54 ;
      RECT 123.18 354.18 123.88 354.34 ;
      RECT 123.18 355.98 123.88 356.14 ;
      RECT 123.24 355.78 123.6 356.14 ;
      RECT 123.24 357.58 123.6 357.94 ;
      RECT 123.18 357.58 123.88 357.74 ;
      RECT 123.18 359.38 123.88 359.54 ;
      RECT 123.24 359.18 123.6 359.54 ;
      RECT 123.24 360.98 123.6 361.34 ;
      RECT 123.18 360.98 123.88 361.14 ;
      RECT 123.18 362.78 123.88 362.94 ;
      RECT 123.24 362.58 123.6 362.94 ;
      RECT 123.24 364.38 123.6 364.74 ;
      RECT 123.18 364.38 123.88 364.54 ;
      RECT 123.18 366.18 123.88 366.34 ;
      RECT 123.24 365.98 123.6 366.34 ;
      RECT 123.24 367.78 123.6 368.14 ;
      RECT 123.18 367.78 123.88 367.94 ;
      RECT 123.18 369.58 123.88 369.74 ;
      RECT 123.24 369.38 123.6 369.74 ;
      RECT 123.24 371.18 123.6 371.54 ;
      RECT 123.18 371.18 123.88 371.34 ;
      RECT 123.18 372.98 123.88 373.14 ;
      RECT 123.24 372.78 123.6 373.14 ;
      RECT 123.24 374.58 123.6 374.94 ;
      RECT 123.18 374.58 123.88 374.74 ;
      RECT 123.18 376.38 123.88 376.54 ;
      RECT 123.24 376.18 123.6 376.54 ;
      RECT 123.24 377.98 123.6 378.34 ;
      RECT 123.18 377.98 123.88 378.14 ;
      RECT 123.18 379.78 123.88 379.94 ;
      RECT 123.24 379.58 123.6 379.94 ;
      RECT 123.24 381.38 123.6 381.74 ;
      RECT 123.18 381.38 123.88 381.54 ;
      RECT 123.18 383.18 123.88 383.34 ;
      RECT 123.24 382.98 123.6 383.34 ;
      RECT 123.24 384.78 123.6 385.14 ;
      RECT 123.18 384.78 123.88 384.94 ;
      RECT 123.18 386.58 123.88 386.74 ;
      RECT 123.24 386.38 123.6 386.74 ;
      RECT 123.24 388.18 123.6 388.54 ;
      RECT 123.18 388.18 123.88 388.34 ;
      RECT 123.18 389.98 123.88 390.14 ;
      RECT 123.24 389.78 123.6 390.14 ;
      RECT 123.24 391.58 123.6 391.94 ;
      RECT 123.18 391.58 123.88 391.74 ;
      RECT 123.18 393.38 123.88 393.54 ;
      RECT 123.24 393.18 123.6 393.54 ;
      RECT 123.24 394.98 123.6 395.34 ;
      RECT 123.18 394.98 123.88 395.14 ;
      RECT 123.18 396.78 123.88 396.94 ;
      RECT 123.24 396.58 123.6 396.94 ;
      RECT 123.24 398.38 123.6 398.74 ;
      RECT 123.18 398.38 123.88 398.54 ;
      RECT 123.18 400.18 123.88 400.34 ;
      RECT 123.24 399.98 123.6 400.34 ;
      RECT 123.24 401.78 123.6 402.14 ;
      RECT 123.18 401.78 123.88 401.94 ;
      RECT 123.18 403.58 123.88 403.74 ;
      RECT 123.24 403.38 123.6 403.74 ;
      RECT 123.24 405.18 123.6 405.54 ;
      RECT 123.18 405.18 123.88 405.34 ;
      RECT 123.18 406.98 123.88 407.14 ;
      RECT 123.24 406.78 123.6 407.14 ;
      RECT 123.24 408.58 123.6 408.94 ;
      RECT 123.18 408.58 123.88 408.74 ;
      RECT 123.18 410.38 123.88 410.54 ;
      RECT 123.24 410.18 123.6 410.54 ;
      RECT 123.24 411.98 123.6 412.34 ;
      RECT 123.18 411.98 123.88 412.14 ;
      RECT 123.18 413.78 123.88 413.94 ;
      RECT 123.24 413.58 123.6 413.94 ;
      RECT 123.24 415.38 123.6 415.74 ;
      RECT 123.18 415.38 123.88 415.54 ;
      RECT 123.18 417.18 123.88 417.34 ;
      RECT 123.24 416.98 123.6 417.34 ;
      RECT 123.24 418.78 123.6 419.14 ;
      RECT 123.18 418.78 123.88 418.94 ;
      RECT 123.18 420.58 123.88 420.74 ;
      RECT 123.24 420.38 123.6 420.74 ;
      RECT 123.24 422.18 123.6 422.54 ;
      RECT 123.18 422.18 123.88 422.34 ;
      RECT 123.18 423.98 123.88 424.14 ;
      RECT 123.24 423.78 123.6 424.14 ;
      RECT 123.24 425.58 123.6 425.94 ;
      RECT 123.18 425.58 123.88 425.74 ;
      RECT 123.18 427.38 123.88 427.54 ;
      RECT 123.24 427.18 123.6 427.54 ;
      RECT 123.24 428.98 123.6 429.34 ;
      RECT 123.18 428.98 123.88 429.14 ;
      RECT 123.18 430.78 123.88 430.94 ;
      RECT 123.24 430.58 123.6 430.94 ;
      RECT 123.24 432.38 123.6 432.74 ;
      RECT 123.18 432.38 123.88 432.54 ;
      RECT 123.18 434.18 123.88 434.34 ;
      RECT 123.24 433.98 123.6 434.34 ;
      RECT 123.24 435.78 123.6 436.14 ;
      RECT 123.18 435.78 123.88 435.94 ;
      RECT 123.18 437.58 123.88 437.74 ;
      RECT 123.24 437.38 123.6 437.74 ;
      RECT 123.24 439.18 123.6 439.54 ;
      RECT 123.18 439.18 123.88 439.34 ;
      RECT 123.18 440.98 123.88 441.14 ;
      RECT 123.24 440.78 123.6 441.14 ;
      RECT 123.24 442.58 123.6 442.94 ;
      RECT 123.18 442.58 123.88 442.74 ;
      RECT 123.18 444.38 123.88 444.54 ;
      RECT 123.24 444.18 123.6 444.54 ;
      RECT 123.24 445.98 123.6 446.34 ;
      RECT 123.18 445.98 123.88 446.14 ;
      RECT 123.18 447.78 123.88 447.94 ;
      RECT 123.24 447.58 123.6 447.94 ;
      RECT 123.24 449.38 123.6 449.74 ;
      RECT 123.18 449.38 123.88 449.54 ;
      RECT 123.18 451.18 123.88 451.34 ;
      RECT 123.24 450.98 123.6 451.34 ;
      RECT 123.24 452.78 123.6 453.14 ;
      RECT 123.18 452.78 123.88 452.94 ;
      RECT 123.18 454.58 123.88 454.74 ;
      RECT 123.24 454.38 123.6 454.74 ;
      RECT 123.24 456.18 123.6 456.54 ;
      RECT 123.18 456.18 123.88 456.34 ;
      RECT 123.18 457.98 123.88 458.14 ;
      RECT 123.24 457.78 123.6 458.14 ;
      RECT 123.24 459.58 123.6 459.94 ;
      RECT 123.18 459.58 123.88 459.74 ;
      RECT 123.18 461.38 123.88 461.54 ;
      RECT 123.24 461.18 123.6 461.54 ;
      RECT 123.24 462.98 123.6 463.34 ;
      RECT 123.18 462.98 123.88 463.14 ;
      RECT 123.18 464.78 123.88 464.94 ;
      RECT 123.24 464.58 123.6 464.94 ;
      RECT 123.24 466.38 123.6 466.74 ;
      RECT 123.18 466.38 123.88 466.54 ;
      RECT 123.18 468.18 123.88 468.34 ;
      RECT 123.24 467.98 123.6 468.34 ;
      RECT 123.24 469.78 123.6 470.14 ;
      RECT 123.18 469.78 123.88 469.94 ;
      RECT 123.18 471.58 123.88 471.74 ;
      RECT 123.24 471.38 123.6 471.74 ;
      RECT 123.24 473.18 123.6 473.54 ;
      RECT 123.18 473.18 123.88 473.34 ;
      RECT 123.18 474.98 123.88 475.14 ;
      RECT 123.24 474.78 123.6 475.14 ;
      RECT 123.24 476.58 123.6 476.94 ;
      RECT 123.18 476.58 123.88 476.74 ;
      RECT 123.18 478.38 123.88 478.54 ;
      RECT 123.24 478.18 123.6 478.54 ;
      RECT 123.24 479.98 123.6 480.34 ;
      RECT 123.18 479.98 123.88 480.14 ;
      RECT 123.18 481.78 123.88 481.94 ;
      RECT 123.24 481.58 123.6 481.94 ;
      RECT 123.24 483.38 123.6 483.74 ;
      RECT 123.18 483.38 123.88 483.54 ;
      RECT 123.18 485.18 123.88 485.34 ;
      RECT 123.24 484.98 123.6 485.34 ;
      RECT 123.24 486.78 123.6 487.14 ;
      RECT 123.18 486.78 123.88 486.94 ;
      RECT 123.18 488.58 123.88 488.74 ;
      RECT 123.24 488.38 123.6 488.74 ;
      RECT 123.24 490.18 123.6 490.54 ;
      RECT 123.18 490.18 123.88 490.34 ;
      RECT 123.18 491.98 123.88 492.14 ;
      RECT 123.24 491.78 123.6 492.14 ;
      RECT 123.24 493.58 123.6 493.94 ;
      RECT 123.18 493.58 123.88 493.74 ;
      RECT 123.18 495.38 123.88 495.54 ;
      RECT 123.24 495.18 123.6 495.54 ;
      RECT 123.24 496.98 123.6 497.34 ;
      RECT 123.18 496.98 123.88 497.14 ;
      RECT 123.18 498.78 123.88 498.94 ;
      RECT 123.24 498.58 123.6 498.94 ;
      RECT 123.24 500.38 123.6 500.74 ;
      RECT 123.18 500.38 123.88 500.54 ;
      RECT 123.18 502.18 123.88 502.34 ;
      RECT 123.24 501.98 123.6 502.34 ;
      RECT 123.24 503.78 123.6 504.14 ;
      RECT 123.18 503.78 123.88 503.94 ;
      RECT 123.55 41.08 123.71 45.17 ;
      RECT 123.55 41.08 123.87 41.24 ;
      RECT 122.55 505.78 123.6 505.94 ;
      RECT 123 505.54 123.6 505.94 ;
      RECT 122.73 31.49 122.89 32.02 ;
      RECT 122.27 31.49 123.35 31.65 ;
      RECT 123.19 27.38 123.35 31.65 ;
      RECT 122.27 27.38 122.43 31.65 ;
      RECT 122.27 27.38 123.35 27.54 ;
      RECT 122.73 26.91 122.89 27.54 ;
      RECT 122.27 51.06 123.35 55.29 ;
      RECT 122.73 50.27 122.89 55.29 ;
      RECT 123.09 49.92 123.25 50.9 ;
      RECT 122.37 49.92 122.53 50.9 ;
      RECT 122.37 49.92 123.25 50.08 ;
      RECT 122.73 45.65 122.89 50.08 ;
      RECT 119.72 72.4 120.72 72.56 ;
      RECT 120.56 71.44 120.72 72.56 ;
      RECT 116.78 72.35 117.66 72.51 ;
      RECT 117.5 71.63 117.66 72.51 ;
      RECT 120.56 72.08 122.97 72.24 ;
      RECT 117.5 71.63 119.24 71.79 ;
      RECT 119.08 71.44 119.24 71.79 ;
      RECT 119.08 71.44 120.72 71.6 ;
      RECT 119.08 74.32 120.72 74.48 ;
      RECT 120.56 73.36 120.72 74.48 ;
      RECT 119.08 74.13 119.24 74.48 ;
      RECT 117.5 74.13 119.24 74.29 ;
      RECT 117.5 73.41 117.66 74.29 ;
      RECT 120.56 73.68 122.97 73.84 ;
      RECT 116.78 73.41 117.66 73.57 ;
      RECT 119.72 73.36 120.72 73.52 ;
      RECT 119.72 79.2 120.72 79.36 ;
      RECT 120.56 78.24 120.72 79.36 ;
      RECT 116.78 79.15 117.66 79.31 ;
      RECT 117.5 78.43 117.66 79.31 ;
      RECT 120.56 78.88 122.97 79.04 ;
      RECT 117.5 78.43 119.24 78.59 ;
      RECT 119.08 78.24 119.24 78.59 ;
      RECT 119.08 78.24 120.72 78.4 ;
      RECT 119.08 81.12 120.72 81.28 ;
      RECT 120.56 80.16 120.72 81.28 ;
      RECT 119.08 80.93 119.24 81.28 ;
      RECT 117.5 80.93 119.24 81.09 ;
      RECT 117.5 80.21 117.66 81.09 ;
      RECT 120.56 80.48 122.97 80.64 ;
      RECT 116.78 80.21 117.66 80.37 ;
      RECT 119.72 80.16 120.72 80.32 ;
      RECT 119.72 86 120.72 86.16 ;
      RECT 120.56 85.04 120.72 86.16 ;
      RECT 116.78 85.95 117.66 86.11 ;
      RECT 117.5 85.23 117.66 86.11 ;
      RECT 120.56 85.68 122.97 85.84 ;
      RECT 117.5 85.23 119.24 85.39 ;
      RECT 119.08 85.04 119.24 85.39 ;
      RECT 119.08 85.04 120.72 85.2 ;
      RECT 119.08 87.92 120.72 88.08 ;
      RECT 120.56 86.96 120.72 88.08 ;
      RECT 119.08 87.73 119.24 88.08 ;
      RECT 117.5 87.73 119.24 87.89 ;
      RECT 117.5 87.01 117.66 87.89 ;
      RECT 120.56 87.28 122.97 87.44 ;
      RECT 116.78 87.01 117.66 87.17 ;
      RECT 119.72 86.96 120.72 87.12 ;
      RECT 119.72 92.8 120.72 92.96 ;
      RECT 120.56 91.84 120.72 92.96 ;
      RECT 116.78 92.75 117.66 92.91 ;
      RECT 117.5 92.03 117.66 92.91 ;
      RECT 120.56 92.48 122.97 92.64 ;
      RECT 117.5 92.03 119.24 92.19 ;
      RECT 119.08 91.84 119.24 92.19 ;
      RECT 119.08 91.84 120.72 92 ;
      RECT 119.08 94.72 120.72 94.88 ;
      RECT 120.56 93.76 120.72 94.88 ;
      RECT 119.08 94.53 119.24 94.88 ;
      RECT 117.5 94.53 119.24 94.69 ;
      RECT 117.5 93.81 117.66 94.69 ;
      RECT 120.56 94.08 122.97 94.24 ;
      RECT 116.78 93.81 117.66 93.97 ;
      RECT 119.72 93.76 120.72 93.92 ;
      RECT 119.72 99.6 120.72 99.76 ;
      RECT 120.56 98.64 120.72 99.76 ;
      RECT 116.78 99.55 117.66 99.71 ;
      RECT 117.5 98.83 117.66 99.71 ;
      RECT 120.56 99.28 122.97 99.44 ;
      RECT 117.5 98.83 119.24 98.99 ;
      RECT 119.08 98.64 119.24 98.99 ;
      RECT 119.08 98.64 120.72 98.8 ;
      RECT 119.08 101.52 120.72 101.68 ;
      RECT 120.56 100.56 120.72 101.68 ;
      RECT 119.08 101.33 119.24 101.68 ;
      RECT 117.5 101.33 119.24 101.49 ;
      RECT 117.5 100.61 117.66 101.49 ;
      RECT 120.56 100.88 122.97 101.04 ;
      RECT 116.78 100.61 117.66 100.77 ;
      RECT 119.72 100.56 120.72 100.72 ;
      RECT 119.72 106.4 120.72 106.56 ;
      RECT 120.56 105.44 120.72 106.56 ;
      RECT 116.78 106.35 117.66 106.51 ;
      RECT 117.5 105.63 117.66 106.51 ;
      RECT 120.56 106.08 122.97 106.24 ;
      RECT 117.5 105.63 119.24 105.79 ;
      RECT 119.08 105.44 119.24 105.79 ;
      RECT 119.08 105.44 120.72 105.6 ;
      RECT 119.08 108.32 120.72 108.48 ;
      RECT 120.56 107.36 120.72 108.48 ;
      RECT 119.08 108.13 119.24 108.48 ;
      RECT 117.5 108.13 119.24 108.29 ;
      RECT 117.5 107.41 117.66 108.29 ;
      RECT 120.56 107.68 122.97 107.84 ;
      RECT 116.78 107.41 117.66 107.57 ;
      RECT 119.72 107.36 120.72 107.52 ;
      RECT 119.72 113.2 120.72 113.36 ;
      RECT 120.56 112.24 120.72 113.36 ;
      RECT 116.78 113.15 117.66 113.31 ;
      RECT 117.5 112.43 117.66 113.31 ;
      RECT 120.56 112.88 122.97 113.04 ;
      RECT 117.5 112.43 119.24 112.59 ;
      RECT 119.08 112.24 119.24 112.59 ;
      RECT 119.08 112.24 120.72 112.4 ;
      RECT 119.08 115.12 120.72 115.28 ;
      RECT 120.56 114.16 120.72 115.28 ;
      RECT 119.08 114.93 119.24 115.28 ;
      RECT 117.5 114.93 119.24 115.09 ;
      RECT 117.5 114.21 117.66 115.09 ;
      RECT 120.56 114.48 122.97 114.64 ;
      RECT 116.78 114.21 117.66 114.37 ;
      RECT 119.72 114.16 120.72 114.32 ;
      RECT 119.72 120 120.72 120.16 ;
      RECT 120.56 119.04 120.72 120.16 ;
      RECT 116.78 119.95 117.66 120.11 ;
      RECT 117.5 119.23 117.66 120.11 ;
      RECT 120.56 119.68 122.97 119.84 ;
      RECT 117.5 119.23 119.24 119.39 ;
      RECT 119.08 119.04 119.24 119.39 ;
      RECT 119.08 119.04 120.72 119.2 ;
      RECT 119.08 121.92 120.72 122.08 ;
      RECT 120.56 120.96 120.72 122.08 ;
      RECT 119.08 121.73 119.24 122.08 ;
      RECT 117.5 121.73 119.24 121.89 ;
      RECT 117.5 121.01 117.66 121.89 ;
      RECT 120.56 121.28 122.97 121.44 ;
      RECT 116.78 121.01 117.66 121.17 ;
      RECT 119.72 120.96 120.72 121.12 ;
      RECT 119.72 126.8 120.72 126.96 ;
      RECT 120.56 125.84 120.72 126.96 ;
      RECT 116.78 126.75 117.66 126.91 ;
      RECT 117.5 126.03 117.66 126.91 ;
      RECT 120.56 126.48 122.97 126.64 ;
      RECT 117.5 126.03 119.24 126.19 ;
      RECT 119.08 125.84 119.24 126.19 ;
      RECT 119.08 125.84 120.72 126 ;
      RECT 119.08 128.72 120.72 128.88 ;
      RECT 120.56 127.76 120.72 128.88 ;
      RECT 119.08 128.53 119.24 128.88 ;
      RECT 117.5 128.53 119.24 128.69 ;
      RECT 117.5 127.81 117.66 128.69 ;
      RECT 120.56 128.08 122.97 128.24 ;
      RECT 116.78 127.81 117.66 127.97 ;
      RECT 119.72 127.76 120.72 127.92 ;
      RECT 119.72 133.6 120.72 133.76 ;
      RECT 120.56 132.64 120.72 133.76 ;
      RECT 116.78 133.55 117.66 133.71 ;
      RECT 117.5 132.83 117.66 133.71 ;
      RECT 120.56 133.28 122.97 133.44 ;
      RECT 117.5 132.83 119.24 132.99 ;
      RECT 119.08 132.64 119.24 132.99 ;
      RECT 119.08 132.64 120.72 132.8 ;
      RECT 119.08 135.52 120.72 135.68 ;
      RECT 120.56 134.56 120.72 135.68 ;
      RECT 119.08 135.33 119.24 135.68 ;
      RECT 117.5 135.33 119.24 135.49 ;
      RECT 117.5 134.61 117.66 135.49 ;
      RECT 120.56 134.88 122.97 135.04 ;
      RECT 116.78 134.61 117.66 134.77 ;
      RECT 119.72 134.56 120.72 134.72 ;
      RECT 119.72 140.4 120.72 140.56 ;
      RECT 120.56 139.44 120.72 140.56 ;
      RECT 116.78 140.35 117.66 140.51 ;
      RECT 117.5 139.63 117.66 140.51 ;
      RECT 120.56 140.08 122.97 140.24 ;
      RECT 117.5 139.63 119.24 139.79 ;
      RECT 119.08 139.44 119.24 139.79 ;
      RECT 119.08 139.44 120.72 139.6 ;
      RECT 119.08 142.32 120.72 142.48 ;
      RECT 120.56 141.36 120.72 142.48 ;
      RECT 119.08 142.13 119.24 142.48 ;
      RECT 117.5 142.13 119.24 142.29 ;
      RECT 117.5 141.41 117.66 142.29 ;
      RECT 120.56 141.68 122.97 141.84 ;
      RECT 116.78 141.41 117.66 141.57 ;
      RECT 119.72 141.36 120.72 141.52 ;
      RECT 119.72 147.2 120.72 147.36 ;
      RECT 120.56 146.24 120.72 147.36 ;
      RECT 116.78 147.15 117.66 147.31 ;
      RECT 117.5 146.43 117.66 147.31 ;
      RECT 120.56 146.88 122.97 147.04 ;
      RECT 117.5 146.43 119.24 146.59 ;
      RECT 119.08 146.24 119.24 146.59 ;
      RECT 119.08 146.24 120.72 146.4 ;
      RECT 119.08 149.12 120.72 149.28 ;
      RECT 120.56 148.16 120.72 149.28 ;
      RECT 119.08 148.93 119.24 149.28 ;
      RECT 117.5 148.93 119.24 149.09 ;
      RECT 117.5 148.21 117.66 149.09 ;
      RECT 120.56 148.48 122.97 148.64 ;
      RECT 116.78 148.21 117.66 148.37 ;
      RECT 119.72 148.16 120.72 148.32 ;
      RECT 119.72 154 120.72 154.16 ;
      RECT 120.56 153.04 120.72 154.16 ;
      RECT 116.78 153.95 117.66 154.11 ;
      RECT 117.5 153.23 117.66 154.11 ;
      RECT 120.56 153.68 122.97 153.84 ;
      RECT 117.5 153.23 119.24 153.39 ;
      RECT 119.08 153.04 119.24 153.39 ;
      RECT 119.08 153.04 120.72 153.2 ;
      RECT 119.08 155.92 120.72 156.08 ;
      RECT 120.56 154.96 120.72 156.08 ;
      RECT 119.08 155.73 119.24 156.08 ;
      RECT 117.5 155.73 119.24 155.89 ;
      RECT 117.5 155.01 117.66 155.89 ;
      RECT 120.56 155.28 122.97 155.44 ;
      RECT 116.78 155.01 117.66 155.17 ;
      RECT 119.72 154.96 120.72 155.12 ;
      RECT 119.72 160.8 120.72 160.96 ;
      RECT 120.56 159.84 120.72 160.96 ;
      RECT 116.78 160.75 117.66 160.91 ;
      RECT 117.5 160.03 117.66 160.91 ;
      RECT 120.56 160.48 122.97 160.64 ;
      RECT 117.5 160.03 119.24 160.19 ;
      RECT 119.08 159.84 119.24 160.19 ;
      RECT 119.08 159.84 120.72 160 ;
      RECT 119.08 162.72 120.72 162.88 ;
      RECT 120.56 161.76 120.72 162.88 ;
      RECT 119.08 162.53 119.24 162.88 ;
      RECT 117.5 162.53 119.24 162.69 ;
      RECT 117.5 161.81 117.66 162.69 ;
      RECT 120.56 162.08 122.97 162.24 ;
      RECT 116.78 161.81 117.66 161.97 ;
      RECT 119.72 161.76 120.72 161.92 ;
      RECT 119.72 167.6 120.72 167.76 ;
      RECT 120.56 166.64 120.72 167.76 ;
      RECT 116.78 167.55 117.66 167.71 ;
      RECT 117.5 166.83 117.66 167.71 ;
      RECT 120.56 167.28 122.97 167.44 ;
      RECT 117.5 166.83 119.24 166.99 ;
      RECT 119.08 166.64 119.24 166.99 ;
      RECT 119.08 166.64 120.72 166.8 ;
      RECT 119.08 169.52 120.72 169.68 ;
      RECT 120.56 168.56 120.72 169.68 ;
      RECT 119.08 169.33 119.24 169.68 ;
      RECT 117.5 169.33 119.24 169.49 ;
      RECT 117.5 168.61 117.66 169.49 ;
      RECT 120.56 168.88 122.97 169.04 ;
      RECT 116.78 168.61 117.66 168.77 ;
      RECT 119.72 168.56 120.72 168.72 ;
      RECT 119.72 174.4 120.72 174.56 ;
      RECT 120.56 173.44 120.72 174.56 ;
      RECT 116.78 174.35 117.66 174.51 ;
      RECT 117.5 173.63 117.66 174.51 ;
      RECT 120.56 174.08 122.97 174.24 ;
      RECT 117.5 173.63 119.24 173.79 ;
      RECT 119.08 173.44 119.24 173.79 ;
      RECT 119.08 173.44 120.72 173.6 ;
      RECT 119.08 176.32 120.72 176.48 ;
      RECT 120.56 175.36 120.72 176.48 ;
      RECT 119.08 176.13 119.24 176.48 ;
      RECT 117.5 176.13 119.24 176.29 ;
      RECT 117.5 175.41 117.66 176.29 ;
      RECT 120.56 175.68 122.97 175.84 ;
      RECT 116.78 175.41 117.66 175.57 ;
      RECT 119.72 175.36 120.72 175.52 ;
      RECT 119.72 181.2 120.72 181.36 ;
      RECT 120.56 180.24 120.72 181.36 ;
      RECT 116.78 181.15 117.66 181.31 ;
      RECT 117.5 180.43 117.66 181.31 ;
      RECT 120.56 180.88 122.97 181.04 ;
      RECT 117.5 180.43 119.24 180.59 ;
      RECT 119.08 180.24 119.24 180.59 ;
      RECT 119.08 180.24 120.72 180.4 ;
      RECT 119.08 183.12 120.72 183.28 ;
      RECT 120.56 182.16 120.72 183.28 ;
      RECT 119.08 182.93 119.24 183.28 ;
      RECT 117.5 182.93 119.24 183.09 ;
      RECT 117.5 182.21 117.66 183.09 ;
      RECT 120.56 182.48 122.97 182.64 ;
      RECT 116.78 182.21 117.66 182.37 ;
      RECT 119.72 182.16 120.72 182.32 ;
      RECT 119.72 188 120.72 188.16 ;
      RECT 120.56 187.04 120.72 188.16 ;
      RECT 116.78 187.95 117.66 188.11 ;
      RECT 117.5 187.23 117.66 188.11 ;
      RECT 120.56 187.68 122.97 187.84 ;
      RECT 117.5 187.23 119.24 187.39 ;
      RECT 119.08 187.04 119.24 187.39 ;
      RECT 119.08 187.04 120.72 187.2 ;
      RECT 119.08 189.92 120.72 190.08 ;
      RECT 120.56 188.96 120.72 190.08 ;
      RECT 119.08 189.73 119.24 190.08 ;
      RECT 117.5 189.73 119.24 189.89 ;
      RECT 117.5 189.01 117.66 189.89 ;
      RECT 120.56 189.28 122.97 189.44 ;
      RECT 116.78 189.01 117.66 189.17 ;
      RECT 119.72 188.96 120.72 189.12 ;
      RECT 119.72 194.8 120.72 194.96 ;
      RECT 120.56 193.84 120.72 194.96 ;
      RECT 116.78 194.75 117.66 194.91 ;
      RECT 117.5 194.03 117.66 194.91 ;
      RECT 120.56 194.48 122.97 194.64 ;
      RECT 117.5 194.03 119.24 194.19 ;
      RECT 119.08 193.84 119.24 194.19 ;
      RECT 119.08 193.84 120.72 194 ;
      RECT 119.08 196.72 120.72 196.88 ;
      RECT 120.56 195.76 120.72 196.88 ;
      RECT 119.08 196.53 119.24 196.88 ;
      RECT 117.5 196.53 119.24 196.69 ;
      RECT 117.5 195.81 117.66 196.69 ;
      RECT 120.56 196.08 122.97 196.24 ;
      RECT 116.78 195.81 117.66 195.97 ;
      RECT 119.72 195.76 120.72 195.92 ;
      RECT 119.72 201.6 120.72 201.76 ;
      RECT 120.56 200.64 120.72 201.76 ;
      RECT 116.78 201.55 117.66 201.71 ;
      RECT 117.5 200.83 117.66 201.71 ;
      RECT 120.56 201.28 122.97 201.44 ;
      RECT 117.5 200.83 119.24 200.99 ;
      RECT 119.08 200.64 119.24 200.99 ;
      RECT 119.08 200.64 120.72 200.8 ;
      RECT 119.08 203.52 120.72 203.68 ;
      RECT 120.56 202.56 120.72 203.68 ;
      RECT 119.08 203.33 119.24 203.68 ;
      RECT 117.5 203.33 119.24 203.49 ;
      RECT 117.5 202.61 117.66 203.49 ;
      RECT 120.56 202.88 122.97 203.04 ;
      RECT 116.78 202.61 117.66 202.77 ;
      RECT 119.72 202.56 120.72 202.72 ;
      RECT 119.72 208.4 120.72 208.56 ;
      RECT 120.56 207.44 120.72 208.56 ;
      RECT 116.78 208.35 117.66 208.51 ;
      RECT 117.5 207.63 117.66 208.51 ;
      RECT 120.56 208.08 122.97 208.24 ;
      RECT 117.5 207.63 119.24 207.79 ;
      RECT 119.08 207.44 119.24 207.79 ;
      RECT 119.08 207.44 120.72 207.6 ;
      RECT 119.08 210.32 120.72 210.48 ;
      RECT 120.56 209.36 120.72 210.48 ;
      RECT 119.08 210.13 119.24 210.48 ;
      RECT 117.5 210.13 119.24 210.29 ;
      RECT 117.5 209.41 117.66 210.29 ;
      RECT 120.56 209.68 122.97 209.84 ;
      RECT 116.78 209.41 117.66 209.57 ;
      RECT 119.72 209.36 120.72 209.52 ;
      RECT 119.72 215.2 120.72 215.36 ;
      RECT 120.56 214.24 120.72 215.36 ;
      RECT 116.78 215.15 117.66 215.31 ;
      RECT 117.5 214.43 117.66 215.31 ;
      RECT 120.56 214.88 122.97 215.04 ;
      RECT 117.5 214.43 119.24 214.59 ;
      RECT 119.08 214.24 119.24 214.59 ;
      RECT 119.08 214.24 120.72 214.4 ;
      RECT 119.08 217.12 120.72 217.28 ;
      RECT 120.56 216.16 120.72 217.28 ;
      RECT 119.08 216.93 119.24 217.28 ;
      RECT 117.5 216.93 119.24 217.09 ;
      RECT 117.5 216.21 117.66 217.09 ;
      RECT 120.56 216.48 122.97 216.64 ;
      RECT 116.78 216.21 117.66 216.37 ;
      RECT 119.72 216.16 120.72 216.32 ;
      RECT 119.72 222 120.72 222.16 ;
      RECT 120.56 221.04 120.72 222.16 ;
      RECT 116.78 221.95 117.66 222.11 ;
      RECT 117.5 221.23 117.66 222.11 ;
      RECT 120.56 221.68 122.97 221.84 ;
      RECT 117.5 221.23 119.24 221.39 ;
      RECT 119.08 221.04 119.24 221.39 ;
      RECT 119.08 221.04 120.72 221.2 ;
      RECT 119.08 223.92 120.72 224.08 ;
      RECT 120.56 222.96 120.72 224.08 ;
      RECT 119.08 223.73 119.24 224.08 ;
      RECT 117.5 223.73 119.24 223.89 ;
      RECT 117.5 223.01 117.66 223.89 ;
      RECT 120.56 223.28 122.97 223.44 ;
      RECT 116.78 223.01 117.66 223.17 ;
      RECT 119.72 222.96 120.72 223.12 ;
      RECT 119.72 228.8 120.72 228.96 ;
      RECT 120.56 227.84 120.72 228.96 ;
      RECT 116.78 228.75 117.66 228.91 ;
      RECT 117.5 228.03 117.66 228.91 ;
      RECT 120.56 228.48 122.97 228.64 ;
      RECT 117.5 228.03 119.24 228.19 ;
      RECT 119.08 227.84 119.24 228.19 ;
      RECT 119.08 227.84 120.72 228 ;
      RECT 119.08 230.72 120.72 230.88 ;
      RECT 120.56 229.76 120.72 230.88 ;
      RECT 119.08 230.53 119.24 230.88 ;
      RECT 117.5 230.53 119.24 230.69 ;
      RECT 117.5 229.81 117.66 230.69 ;
      RECT 120.56 230.08 122.97 230.24 ;
      RECT 116.78 229.81 117.66 229.97 ;
      RECT 119.72 229.76 120.72 229.92 ;
      RECT 119.72 235.6 120.72 235.76 ;
      RECT 120.56 234.64 120.72 235.76 ;
      RECT 116.78 235.55 117.66 235.71 ;
      RECT 117.5 234.83 117.66 235.71 ;
      RECT 120.56 235.28 122.97 235.44 ;
      RECT 117.5 234.83 119.24 234.99 ;
      RECT 119.08 234.64 119.24 234.99 ;
      RECT 119.08 234.64 120.72 234.8 ;
      RECT 119.08 237.52 120.72 237.68 ;
      RECT 120.56 236.56 120.72 237.68 ;
      RECT 119.08 237.33 119.24 237.68 ;
      RECT 117.5 237.33 119.24 237.49 ;
      RECT 117.5 236.61 117.66 237.49 ;
      RECT 120.56 236.88 122.97 237.04 ;
      RECT 116.78 236.61 117.66 236.77 ;
      RECT 119.72 236.56 120.72 236.72 ;
      RECT 119.72 242.4 120.72 242.56 ;
      RECT 120.56 241.44 120.72 242.56 ;
      RECT 116.78 242.35 117.66 242.51 ;
      RECT 117.5 241.63 117.66 242.51 ;
      RECT 120.56 242.08 122.97 242.24 ;
      RECT 117.5 241.63 119.24 241.79 ;
      RECT 119.08 241.44 119.24 241.79 ;
      RECT 119.08 241.44 120.72 241.6 ;
      RECT 119.08 244.32 120.72 244.48 ;
      RECT 120.56 243.36 120.72 244.48 ;
      RECT 119.08 244.13 119.24 244.48 ;
      RECT 117.5 244.13 119.24 244.29 ;
      RECT 117.5 243.41 117.66 244.29 ;
      RECT 120.56 243.68 122.97 243.84 ;
      RECT 116.78 243.41 117.66 243.57 ;
      RECT 119.72 243.36 120.72 243.52 ;
      RECT 119.72 249.2 120.72 249.36 ;
      RECT 120.56 248.24 120.72 249.36 ;
      RECT 116.78 249.15 117.66 249.31 ;
      RECT 117.5 248.43 117.66 249.31 ;
      RECT 120.56 248.88 122.97 249.04 ;
      RECT 117.5 248.43 119.24 248.59 ;
      RECT 119.08 248.24 119.24 248.59 ;
      RECT 119.08 248.24 120.72 248.4 ;
      RECT 119.08 251.12 120.72 251.28 ;
      RECT 120.56 250.16 120.72 251.28 ;
      RECT 119.08 250.93 119.24 251.28 ;
      RECT 117.5 250.93 119.24 251.09 ;
      RECT 117.5 250.21 117.66 251.09 ;
      RECT 120.56 250.48 122.97 250.64 ;
      RECT 116.78 250.21 117.66 250.37 ;
      RECT 119.72 250.16 120.72 250.32 ;
      RECT 119.72 256 120.72 256.16 ;
      RECT 120.56 255.04 120.72 256.16 ;
      RECT 116.78 255.95 117.66 256.11 ;
      RECT 117.5 255.23 117.66 256.11 ;
      RECT 120.56 255.68 122.97 255.84 ;
      RECT 117.5 255.23 119.24 255.39 ;
      RECT 119.08 255.04 119.24 255.39 ;
      RECT 119.08 255.04 120.72 255.2 ;
      RECT 119.08 257.92 120.72 258.08 ;
      RECT 120.56 256.96 120.72 258.08 ;
      RECT 119.08 257.73 119.24 258.08 ;
      RECT 117.5 257.73 119.24 257.89 ;
      RECT 117.5 257.01 117.66 257.89 ;
      RECT 120.56 257.28 122.97 257.44 ;
      RECT 116.78 257.01 117.66 257.17 ;
      RECT 119.72 256.96 120.72 257.12 ;
      RECT 119.72 262.8 120.72 262.96 ;
      RECT 120.56 261.84 120.72 262.96 ;
      RECT 116.78 262.75 117.66 262.91 ;
      RECT 117.5 262.03 117.66 262.91 ;
      RECT 120.56 262.48 122.97 262.64 ;
      RECT 117.5 262.03 119.24 262.19 ;
      RECT 119.08 261.84 119.24 262.19 ;
      RECT 119.08 261.84 120.72 262 ;
      RECT 119.08 264.72 120.72 264.88 ;
      RECT 120.56 263.76 120.72 264.88 ;
      RECT 119.08 264.53 119.24 264.88 ;
      RECT 117.5 264.53 119.24 264.69 ;
      RECT 117.5 263.81 117.66 264.69 ;
      RECT 120.56 264.08 122.97 264.24 ;
      RECT 116.78 263.81 117.66 263.97 ;
      RECT 119.72 263.76 120.72 263.92 ;
      RECT 119.72 269.6 120.72 269.76 ;
      RECT 120.56 268.64 120.72 269.76 ;
      RECT 116.78 269.55 117.66 269.71 ;
      RECT 117.5 268.83 117.66 269.71 ;
      RECT 120.56 269.28 122.97 269.44 ;
      RECT 117.5 268.83 119.24 268.99 ;
      RECT 119.08 268.64 119.24 268.99 ;
      RECT 119.08 268.64 120.72 268.8 ;
      RECT 119.08 271.52 120.72 271.68 ;
      RECT 120.56 270.56 120.72 271.68 ;
      RECT 119.08 271.33 119.24 271.68 ;
      RECT 117.5 271.33 119.24 271.49 ;
      RECT 117.5 270.61 117.66 271.49 ;
      RECT 120.56 270.88 122.97 271.04 ;
      RECT 116.78 270.61 117.66 270.77 ;
      RECT 119.72 270.56 120.72 270.72 ;
      RECT 119.72 276.4 120.72 276.56 ;
      RECT 120.56 275.44 120.72 276.56 ;
      RECT 116.78 276.35 117.66 276.51 ;
      RECT 117.5 275.63 117.66 276.51 ;
      RECT 120.56 276.08 122.97 276.24 ;
      RECT 117.5 275.63 119.24 275.79 ;
      RECT 119.08 275.44 119.24 275.79 ;
      RECT 119.08 275.44 120.72 275.6 ;
      RECT 119.08 278.32 120.72 278.48 ;
      RECT 120.56 277.36 120.72 278.48 ;
      RECT 119.08 278.13 119.24 278.48 ;
      RECT 117.5 278.13 119.24 278.29 ;
      RECT 117.5 277.41 117.66 278.29 ;
      RECT 120.56 277.68 122.97 277.84 ;
      RECT 116.78 277.41 117.66 277.57 ;
      RECT 119.72 277.36 120.72 277.52 ;
      RECT 119.72 283.2 120.72 283.36 ;
      RECT 120.56 282.24 120.72 283.36 ;
      RECT 116.78 283.15 117.66 283.31 ;
      RECT 117.5 282.43 117.66 283.31 ;
      RECT 120.56 282.88 122.97 283.04 ;
      RECT 117.5 282.43 119.24 282.59 ;
      RECT 119.08 282.24 119.24 282.59 ;
      RECT 119.08 282.24 120.72 282.4 ;
      RECT 119.08 285.12 120.72 285.28 ;
      RECT 120.56 284.16 120.72 285.28 ;
      RECT 119.08 284.93 119.24 285.28 ;
      RECT 117.5 284.93 119.24 285.09 ;
      RECT 117.5 284.21 117.66 285.09 ;
      RECT 120.56 284.48 122.97 284.64 ;
      RECT 116.78 284.21 117.66 284.37 ;
      RECT 119.72 284.16 120.72 284.32 ;
      RECT 119.72 290 120.72 290.16 ;
      RECT 120.56 289.04 120.72 290.16 ;
      RECT 116.78 289.95 117.66 290.11 ;
      RECT 117.5 289.23 117.66 290.11 ;
      RECT 120.56 289.68 122.97 289.84 ;
      RECT 117.5 289.23 119.24 289.39 ;
      RECT 119.08 289.04 119.24 289.39 ;
      RECT 119.08 289.04 120.72 289.2 ;
      RECT 119.08 291.92 120.72 292.08 ;
      RECT 120.56 290.96 120.72 292.08 ;
      RECT 119.08 291.73 119.24 292.08 ;
      RECT 117.5 291.73 119.24 291.89 ;
      RECT 117.5 291.01 117.66 291.89 ;
      RECT 120.56 291.28 122.97 291.44 ;
      RECT 116.78 291.01 117.66 291.17 ;
      RECT 119.72 290.96 120.72 291.12 ;
      RECT 119.72 296.8 120.72 296.96 ;
      RECT 120.56 295.84 120.72 296.96 ;
      RECT 116.78 296.75 117.66 296.91 ;
      RECT 117.5 296.03 117.66 296.91 ;
      RECT 120.56 296.48 122.97 296.64 ;
      RECT 117.5 296.03 119.24 296.19 ;
      RECT 119.08 295.84 119.24 296.19 ;
      RECT 119.08 295.84 120.72 296 ;
      RECT 119.08 298.72 120.72 298.88 ;
      RECT 120.56 297.76 120.72 298.88 ;
      RECT 119.08 298.53 119.24 298.88 ;
      RECT 117.5 298.53 119.24 298.69 ;
      RECT 117.5 297.81 117.66 298.69 ;
      RECT 120.56 298.08 122.97 298.24 ;
      RECT 116.78 297.81 117.66 297.97 ;
      RECT 119.72 297.76 120.72 297.92 ;
      RECT 119.72 303.6 120.72 303.76 ;
      RECT 120.56 302.64 120.72 303.76 ;
      RECT 116.78 303.55 117.66 303.71 ;
      RECT 117.5 302.83 117.66 303.71 ;
      RECT 120.56 303.28 122.97 303.44 ;
      RECT 117.5 302.83 119.24 302.99 ;
      RECT 119.08 302.64 119.24 302.99 ;
      RECT 119.08 302.64 120.72 302.8 ;
      RECT 119.08 305.52 120.72 305.68 ;
      RECT 120.56 304.56 120.72 305.68 ;
      RECT 119.08 305.33 119.24 305.68 ;
      RECT 117.5 305.33 119.24 305.49 ;
      RECT 117.5 304.61 117.66 305.49 ;
      RECT 120.56 304.88 122.97 305.04 ;
      RECT 116.78 304.61 117.66 304.77 ;
      RECT 119.72 304.56 120.72 304.72 ;
      RECT 119.72 310.4 120.72 310.56 ;
      RECT 120.56 309.44 120.72 310.56 ;
      RECT 116.78 310.35 117.66 310.51 ;
      RECT 117.5 309.63 117.66 310.51 ;
      RECT 120.56 310.08 122.97 310.24 ;
      RECT 117.5 309.63 119.24 309.79 ;
      RECT 119.08 309.44 119.24 309.79 ;
      RECT 119.08 309.44 120.72 309.6 ;
      RECT 119.08 312.32 120.72 312.48 ;
      RECT 120.56 311.36 120.72 312.48 ;
      RECT 119.08 312.13 119.24 312.48 ;
      RECT 117.5 312.13 119.24 312.29 ;
      RECT 117.5 311.41 117.66 312.29 ;
      RECT 120.56 311.68 122.97 311.84 ;
      RECT 116.78 311.41 117.66 311.57 ;
      RECT 119.72 311.36 120.72 311.52 ;
      RECT 119.72 317.2 120.72 317.36 ;
      RECT 120.56 316.24 120.72 317.36 ;
      RECT 116.78 317.15 117.66 317.31 ;
      RECT 117.5 316.43 117.66 317.31 ;
      RECT 120.56 316.88 122.97 317.04 ;
      RECT 117.5 316.43 119.24 316.59 ;
      RECT 119.08 316.24 119.24 316.59 ;
      RECT 119.08 316.24 120.72 316.4 ;
      RECT 119.08 319.12 120.72 319.28 ;
      RECT 120.56 318.16 120.72 319.28 ;
      RECT 119.08 318.93 119.24 319.28 ;
      RECT 117.5 318.93 119.24 319.09 ;
      RECT 117.5 318.21 117.66 319.09 ;
      RECT 120.56 318.48 122.97 318.64 ;
      RECT 116.78 318.21 117.66 318.37 ;
      RECT 119.72 318.16 120.72 318.32 ;
      RECT 119.72 324 120.72 324.16 ;
      RECT 120.56 323.04 120.72 324.16 ;
      RECT 116.78 323.95 117.66 324.11 ;
      RECT 117.5 323.23 117.66 324.11 ;
      RECT 120.56 323.68 122.97 323.84 ;
      RECT 117.5 323.23 119.24 323.39 ;
      RECT 119.08 323.04 119.24 323.39 ;
      RECT 119.08 323.04 120.72 323.2 ;
      RECT 119.08 325.92 120.72 326.08 ;
      RECT 120.56 324.96 120.72 326.08 ;
      RECT 119.08 325.73 119.24 326.08 ;
      RECT 117.5 325.73 119.24 325.89 ;
      RECT 117.5 325.01 117.66 325.89 ;
      RECT 120.56 325.28 122.97 325.44 ;
      RECT 116.78 325.01 117.66 325.17 ;
      RECT 119.72 324.96 120.72 325.12 ;
      RECT 119.72 330.8 120.72 330.96 ;
      RECT 120.56 329.84 120.72 330.96 ;
      RECT 116.78 330.75 117.66 330.91 ;
      RECT 117.5 330.03 117.66 330.91 ;
      RECT 120.56 330.48 122.97 330.64 ;
      RECT 117.5 330.03 119.24 330.19 ;
      RECT 119.08 329.84 119.24 330.19 ;
      RECT 119.08 329.84 120.72 330 ;
      RECT 119.08 332.72 120.72 332.88 ;
      RECT 120.56 331.76 120.72 332.88 ;
      RECT 119.08 332.53 119.24 332.88 ;
      RECT 117.5 332.53 119.24 332.69 ;
      RECT 117.5 331.81 117.66 332.69 ;
      RECT 120.56 332.08 122.97 332.24 ;
      RECT 116.78 331.81 117.66 331.97 ;
      RECT 119.72 331.76 120.72 331.92 ;
      RECT 119.72 337.6 120.72 337.76 ;
      RECT 120.56 336.64 120.72 337.76 ;
      RECT 116.78 337.55 117.66 337.71 ;
      RECT 117.5 336.83 117.66 337.71 ;
      RECT 120.56 337.28 122.97 337.44 ;
      RECT 117.5 336.83 119.24 336.99 ;
      RECT 119.08 336.64 119.24 336.99 ;
      RECT 119.08 336.64 120.72 336.8 ;
      RECT 119.08 339.52 120.72 339.68 ;
      RECT 120.56 338.56 120.72 339.68 ;
      RECT 119.08 339.33 119.24 339.68 ;
      RECT 117.5 339.33 119.24 339.49 ;
      RECT 117.5 338.61 117.66 339.49 ;
      RECT 120.56 338.88 122.97 339.04 ;
      RECT 116.78 338.61 117.66 338.77 ;
      RECT 119.72 338.56 120.72 338.72 ;
      RECT 119.72 344.4 120.72 344.56 ;
      RECT 120.56 343.44 120.72 344.56 ;
      RECT 116.78 344.35 117.66 344.51 ;
      RECT 117.5 343.63 117.66 344.51 ;
      RECT 120.56 344.08 122.97 344.24 ;
      RECT 117.5 343.63 119.24 343.79 ;
      RECT 119.08 343.44 119.24 343.79 ;
      RECT 119.08 343.44 120.72 343.6 ;
      RECT 119.08 346.32 120.72 346.48 ;
      RECT 120.56 345.36 120.72 346.48 ;
      RECT 119.08 346.13 119.24 346.48 ;
      RECT 117.5 346.13 119.24 346.29 ;
      RECT 117.5 345.41 117.66 346.29 ;
      RECT 120.56 345.68 122.97 345.84 ;
      RECT 116.78 345.41 117.66 345.57 ;
      RECT 119.72 345.36 120.72 345.52 ;
      RECT 119.72 351.2 120.72 351.36 ;
      RECT 120.56 350.24 120.72 351.36 ;
      RECT 116.78 351.15 117.66 351.31 ;
      RECT 117.5 350.43 117.66 351.31 ;
      RECT 120.56 350.88 122.97 351.04 ;
      RECT 117.5 350.43 119.24 350.59 ;
      RECT 119.08 350.24 119.24 350.59 ;
      RECT 119.08 350.24 120.72 350.4 ;
      RECT 119.08 353.12 120.72 353.28 ;
      RECT 120.56 352.16 120.72 353.28 ;
      RECT 119.08 352.93 119.24 353.28 ;
      RECT 117.5 352.93 119.24 353.09 ;
      RECT 117.5 352.21 117.66 353.09 ;
      RECT 120.56 352.48 122.97 352.64 ;
      RECT 116.78 352.21 117.66 352.37 ;
      RECT 119.72 352.16 120.72 352.32 ;
      RECT 119.72 358 120.72 358.16 ;
      RECT 120.56 357.04 120.72 358.16 ;
      RECT 116.78 357.95 117.66 358.11 ;
      RECT 117.5 357.23 117.66 358.11 ;
      RECT 120.56 357.68 122.97 357.84 ;
      RECT 117.5 357.23 119.24 357.39 ;
      RECT 119.08 357.04 119.24 357.39 ;
      RECT 119.08 357.04 120.72 357.2 ;
      RECT 119.08 359.92 120.72 360.08 ;
      RECT 120.56 358.96 120.72 360.08 ;
      RECT 119.08 359.73 119.24 360.08 ;
      RECT 117.5 359.73 119.24 359.89 ;
      RECT 117.5 359.01 117.66 359.89 ;
      RECT 120.56 359.28 122.97 359.44 ;
      RECT 116.78 359.01 117.66 359.17 ;
      RECT 119.72 358.96 120.72 359.12 ;
      RECT 119.72 364.8 120.72 364.96 ;
      RECT 120.56 363.84 120.72 364.96 ;
      RECT 116.78 364.75 117.66 364.91 ;
      RECT 117.5 364.03 117.66 364.91 ;
      RECT 120.56 364.48 122.97 364.64 ;
      RECT 117.5 364.03 119.24 364.19 ;
      RECT 119.08 363.84 119.24 364.19 ;
      RECT 119.08 363.84 120.72 364 ;
      RECT 119.08 366.72 120.72 366.88 ;
      RECT 120.56 365.76 120.72 366.88 ;
      RECT 119.08 366.53 119.24 366.88 ;
      RECT 117.5 366.53 119.24 366.69 ;
      RECT 117.5 365.81 117.66 366.69 ;
      RECT 120.56 366.08 122.97 366.24 ;
      RECT 116.78 365.81 117.66 365.97 ;
      RECT 119.72 365.76 120.72 365.92 ;
      RECT 119.72 371.6 120.72 371.76 ;
      RECT 120.56 370.64 120.72 371.76 ;
      RECT 116.78 371.55 117.66 371.71 ;
      RECT 117.5 370.83 117.66 371.71 ;
      RECT 120.56 371.28 122.97 371.44 ;
      RECT 117.5 370.83 119.24 370.99 ;
      RECT 119.08 370.64 119.24 370.99 ;
      RECT 119.08 370.64 120.72 370.8 ;
      RECT 119.08 373.52 120.72 373.68 ;
      RECT 120.56 372.56 120.72 373.68 ;
      RECT 119.08 373.33 119.24 373.68 ;
      RECT 117.5 373.33 119.24 373.49 ;
      RECT 117.5 372.61 117.66 373.49 ;
      RECT 120.56 372.88 122.97 373.04 ;
      RECT 116.78 372.61 117.66 372.77 ;
      RECT 119.72 372.56 120.72 372.72 ;
      RECT 119.72 378.4 120.72 378.56 ;
      RECT 120.56 377.44 120.72 378.56 ;
      RECT 116.78 378.35 117.66 378.51 ;
      RECT 117.5 377.63 117.66 378.51 ;
      RECT 120.56 378.08 122.97 378.24 ;
      RECT 117.5 377.63 119.24 377.79 ;
      RECT 119.08 377.44 119.24 377.79 ;
      RECT 119.08 377.44 120.72 377.6 ;
      RECT 119.08 380.32 120.72 380.48 ;
      RECT 120.56 379.36 120.72 380.48 ;
      RECT 119.08 380.13 119.24 380.48 ;
      RECT 117.5 380.13 119.24 380.29 ;
      RECT 117.5 379.41 117.66 380.29 ;
      RECT 120.56 379.68 122.97 379.84 ;
      RECT 116.78 379.41 117.66 379.57 ;
      RECT 119.72 379.36 120.72 379.52 ;
      RECT 119.72 385.2 120.72 385.36 ;
      RECT 120.56 384.24 120.72 385.36 ;
      RECT 116.78 385.15 117.66 385.31 ;
      RECT 117.5 384.43 117.66 385.31 ;
      RECT 120.56 384.88 122.97 385.04 ;
      RECT 117.5 384.43 119.24 384.59 ;
      RECT 119.08 384.24 119.24 384.59 ;
      RECT 119.08 384.24 120.72 384.4 ;
      RECT 119.08 387.12 120.72 387.28 ;
      RECT 120.56 386.16 120.72 387.28 ;
      RECT 119.08 386.93 119.24 387.28 ;
      RECT 117.5 386.93 119.24 387.09 ;
      RECT 117.5 386.21 117.66 387.09 ;
      RECT 120.56 386.48 122.97 386.64 ;
      RECT 116.78 386.21 117.66 386.37 ;
      RECT 119.72 386.16 120.72 386.32 ;
      RECT 119.72 392 120.72 392.16 ;
      RECT 120.56 391.04 120.72 392.16 ;
      RECT 116.78 391.95 117.66 392.11 ;
      RECT 117.5 391.23 117.66 392.11 ;
      RECT 120.56 391.68 122.97 391.84 ;
      RECT 117.5 391.23 119.24 391.39 ;
      RECT 119.08 391.04 119.24 391.39 ;
      RECT 119.08 391.04 120.72 391.2 ;
      RECT 119.08 393.92 120.72 394.08 ;
      RECT 120.56 392.96 120.72 394.08 ;
      RECT 119.08 393.73 119.24 394.08 ;
      RECT 117.5 393.73 119.24 393.89 ;
      RECT 117.5 393.01 117.66 393.89 ;
      RECT 120.56 393.28 122.97 393.44 ;
      RECT 116.78 393.01 117.66 393.17 ;
      RECT 119.72 392.96 120.72 393.12 ;
      RECT 119.72 398.8 120.72 398.96 ;
      RECT 120.56 397.84 120.72 398.96 ;
      RECT 116.78 398.75 117.66 398.91 ;
      RECT 117.5 398.03 117.66 398.91 ;
      RECT 120.56 398.48 122.97 398.64 ;
      RECT 117.5 398.03 119.24 398.19 ;
      RECT 119.08 397.84 119.24 398.19 ;
      RECT 119.08 397.84 120.72 398 ;
      RECT 119.08 400.72 120.72 400.88 ;
      RECT 120.56 399.76 120.72 400.88 ;
      RECT 119.08 400.53 119.24 400.88 ;
      RECT 117.5 400.53 119.24 400.69 ;
      RECT 117.5 399.81 117.66 400.69 ;
      RECT 120.56 400.08 122.97 400.24 ;
      RECT 116.78 399.81 117.66 399.97 ;
      RECT 119.72 399.76 120.72 399.92 ;
      RECT 119.72 405.6 120.72 405.76 ;
      RECT 120.56 404.64 120.72 405.76 ;
      RECT 116.78 405.55 117.66 405.71 ;
      RECT 117.5 404.83 117.66 405.71 ;
      RECT 120.56 405.28 122.97 405.44 ;
      RECT 117.5 404.83 119.24 404.99 ;
      RECT 119.08 404.64 119.24 404.99 ;
      RECT 119.08 404.64 120.72 404.8 ;
      RECT 119.08 407.52 120.72 407.68 ;
      RECT 120.56 406.56 120.72 407.68 ;
      RECT 119.08 407.33 119.24 407.68 ;
      RECT 117.5 407.33 119.24 407.49 ;
      RECT 117.5 406.61 117.66 407.49 ;
      RECT 120.56 406.88 122.97 407.04 ;
      RECT 116.78 406.61 117.66 406.77 ;
      RECT 119.72 406.56 120.72 406.72 ;
      RECT 119.72 412.4 120.72 412.56 ;
      RECT 120.56 411.44 120.72 412.56 ;
      RECT 116.78 412.35 117.66 412.51 ;
      RECT 117.5 411.63 117.66 412.51 ;
      RECT 120.56 412.08 122.97 412.24 ;
      RECT 117.5 411.63 119.24 411.79 ;
      RECT 119.08 411.44 119.24 411.79 ;
      RECT 119.08 411.44 120.72 411.6 ;
      RECT 119.08 414.32 120.72 414.48 ;
      RECT 120.56 413.36 120.72 414.48 ;
      RECT 119.08 414.13 119.24 414.48 ;
      RECT 117.5 414.13 119.24 414.29 ;
      RECT 117.5 413.41 117.66 414.29 ;
      RECT 120.56 413.68 122.97 413.84 ;
      RECT 116.78 413.41 117.66 413.57 ;
      RECT 119.72 413.36 120.72 413.52 ;
      RECT 119.72 419.2 120.72 419.36 ;
      RECT 120.56 418.24 120.72 419.36 ;
      RECT 116.78 419.15 117.66 419.31 ;
      RECT 117.5 418.43 117.66 419.31 ;
      RECT 120.56 418.88 122.97 419.04 ;
      RECT 117.5 418.43 119.24 418.59 ;
      RECT 119.08 418.24 119.24 418.59 ;
      RECT 119.08 418.24 120.72 418.4 ;
      RECT 119.08 421.12 120.72 421.28 ;
      RECT 120.56 420.16 120.72 421.28 ;
      RECT 119.08 420.93 119.24 421.28 ;
      RECT 117.5 420.93 119.24 421.09 ;
      RECT 117.5 420.21 117.66 421.09 ;
      RECT 120.56 420.48 122.97 420.64 ;
      RECT 116.78 420.21 117.66 420.37 ;
      RECT 119.72 420.16 120.72 420.32 ;
      RECT 119.72 426 120.72 426.16 ;
      RECT 120.56 425.04 120.72 426.16 ;
      RECT 116.78 425.95 117.66 426.11 ;
      RECT 117.5 425.23 117.66 426.11 ;
      RECT 120.56 425.68 122.97 425.84 ;
      RECT 117.5 425.23 119.24 425.39 ;
      RECT 119.08 425.04 119.24 425.39 ;
      RECT 119.08 425.04 120.72 425.2 ;
      RECT 119.08 427.92 120.72 428.08 ;
      RECT 120.56 426.96 120.72 428.08 ;
      RECT 119.08 427.73 119.24 428.08 ;
      RECT 117.5 427.73 119.24 427.89 ;
      RECT 117.5 427.01 117.66 427.89 ;
      RECT 120.56 427.28 122.97 427.44 ;
      RECT 116.78 427.01 117.66 427.17 ;
      RECT 119.72 426.96 120.72 427.12 ;
      RECT 119.72 432.8 120.72 432.96 ;
      RECT 120.56 431.84 120.72 432.96 ;
      RECT 116.78 432.75 117.66 432.91 ;
      RECT 117.5 432.03 117.66 432.91 ;
      RECT 120.56 432.48 122.97 432.64 ;
      RECT 117.5 432.03 119.24 432.19 ;
      RECT 119.08 431.84 119.24 432.19 ;
      RECT 119.08 431.84 120.72 432 ;
      RECT 119.08 434.72 120.72 434.88 ;
      RECT 120.56 433.76 120.72 434.88 ;
      RECT 119.08 434.53 119.24 434.88 ;
      RECT 117.5 434.53 119.24 434.69 ;
      RECT 117.5 433.81 117.66 434.69 ;
      RECT 120.56 434.08 122.97 434.24 ;
      RECT 116.78 433.81 117.66 433.97 ;
      RECT 119.72 433.76 120.72 433.92 ;
      RECT 119.72 439.6 120.72 439.76 ;
      RECT 120.56 438.64 120.72 439.76 ;
      RECT 116.78 439.55 117.66 439.71 ;
      RECT 117.5 438.83 117.66 439.71 ;
      RECT 120.56 439.28 122.97 439.44 ;
      RECT 117.5 438.83 119.24 438.99 ;
      RECT 119.08 438.64 119.24 438.99 ;
      RECT 119.08 438.64 120.72 438.8 ;
      RECT 119.08 441.52 120.72 441.68 ;
      RECT 120.56 440.56 120.72 441.68 ;
      RECT 119.08 441.33 119.24 441.68 ;
      RECT 117.5 441.33 119.24 441.49 ;
      RECT 117.5 440.61 117.66 441.49 ;
      RECT 120.56 440.88 122.97 441.04 ;
      RECT 116.78 440.61 117.66 440.77 ;
      RECT 119.72 440.56 120.72 440.72 ;
      RECT 119.72 446.4 120.72 446.56 ;
      RECT 120.56 445.44 120.72 446.56 ;
      RECT 116.78 446.35 117.66 446.51 ;
      RECT 117.5 445.63 117.66 446.51 ;
      RECT 120.56 446.08 122.97 446.24 ;
      RECT 117.5 445.63 119.24 445.79 ;
      RECT 119.08 445.44 119.24 445.79 ;
      RECT 119.08 445.44 120.72 445.6 ;
      RECT 119.08 448.32 120.72 448.48 ;
      RECT 120.56 447.36 120.72 448.48 ;
      RECT 119.08 448.13 119.24 448.48 ;
      RECT 117.5 448.13 119.24 448.29 ;
      RECT 117.5 447.41 117.66 448.29 ;
      RECT 120.56 447.68 122.97 447.84 ;
      RECT 116.78 447.41 117.66 447.57 ;
      RECT 119.72 447.36 120.72 447.52 ;
      RECT 119.72 453.2 120.72 453.36 ;
      RECT 120.56 452.24 120.72 453.36 ;
      RECT 116.78 453.15 117.66 453.31 ;
      RECT 117.5 452.43 117.66 453.31 ;
      RECT 120.56 452.88 122.97 453.04 ;
      RECT 117.5 452.43 119.24 452.59 ;
      RECT 119.08 452.24 119.24 452.59 ;
      RECT 119.08 452.24 120.72 452.4 ;
      RECT 119.08 455.12 120.72 455.28 ;
      RECT 120.56 454.16 120.72 455.28 ;
      RECT 119.08 454.93 119.24 455.28 ;
      RECT 117.5 454.93 119.24 455.09 ;
      RECT 117.5 454.21 117.66 455.09 ;
      RECT 120.56 454.48 122.97 454.64 ;
      RECT 116.78 454.21 117.66 454.37 ;
      RECT 119.72 454.16 120.72 454.32 ;
      RECT 119.72 460 120.72 460.16 ;
      RECT 120.56 459.04 120.72 460.16 ;
      RECT 116.78 459.95 117.66 460.11 ;
      RECT 117.5 459.23 117.66 460.11 ;
      RECT 120.56 459.68 122.97 459.84 ;
      RECT 117.5 459.23 119.24 459.39 ;
      RECT 119.08 459.04 119.24 459.39 ;
      RECT 119.08 459.04 120.72 459.2 ;
      RECT 119.08 461.92 120.72 462.08 ;
      RECT 120.56 460.96 120.72 462.08 ;
      RECT 119.08 461.73 119.24 462.08 ;
      RECT 117.5 461.73 119.24 461.89 ;
      RECT 117.5 461.01 117.66 461.89 ;
      RECT 120.56 461.28 122.97 461.44 ;
      RECT 116.78 461.01 117.66 461.17 ;
      RECT 119.72 460.96 120.72 461.12 ;
      RECT 119.72 466.8 120.72 466.96 ;
      RECT 120.56 465.84 120.72 466.96 ;
      RECT 116.78 466.75 117.66 466.91 ;
      RECT 117.5 466.03 117.66 466.91 ;
      RECT 120.56 466.48 122.97 466.64 ;
      RECT 117.5 466.03 119.24 466.19 ;
      RECT 119.08 465.84 119.24 466.19 ;
      RECT 119.08 465.84 120.72 466 ;
      RECT 119.08 468.72 120.72 468.88 ;
      RECT 120.56 467.76 120.72 468.88 ;
      RECT 119.08 468.53 119.24 468.88 ;
      RECT 117.5 468.53 119.24 468.69 ;
      RECT 117.5 467.81 117.66 468.69 ;
      RECT 120.56 468.08 122.97 468.24 ;
      RECT 116.78 467.81 117.66 467.97 ;
      RECT 119.72 467.76 120.72 467.92 ;
      RECT 119.72 473.6 120.72 473.76 ;
      RECT 120.56 472.64 120.72 473.76 ;
      RECT 116.78 473.55 117.66 473.71 ;
      RECT 117.5 472.83 117.66 473.71 ;
      RECT 120.56 473.28 122.97 473.44 ;
      RECT 117.5 472.83 119.24 472.99 ;
      RECT 119.08 472.64 119.24 472.99 ;
      RECT 119.08 472.64 120.72 472.8 ;
      RECT 119.08 475.52 120.72 475.68 ;
      RECT 120.56 474.56 120.72 475.68 ;
      RECT 119.08 475.33 119.24 475.68 ;
      RECT 117.5 475.33 119.24 475.49 ;
      RECT 117.5 474.61 117.66 475.49 ;
      RECT 120.56 474.88 122.97 475.04 ;
      RECT 116.78 474.61 117.66 474.77 ;
      RECT 119.72 474.56 120.72 474.72 ;
      RECT 119.72 480.4 120.72 480.56 ;
      RECT 120.56 479.44 120.72 480.56 ;
      RECT 116.78 480.35 117.66 480.51 ;
      RECT 117.5 479.63 117.66 480.51 ;
      RECT 120.56 480.08 122.97 480.24 ;
      RECT 117.5 479.63 119.24 479.79 ;
      RECT 119.08 479.44 119.24 479.79 ;
      RECT 119.08 479.44 120.72 479.6 ;
      RECT 119.08 482.32 120.72 482.48 ;
      RECT 120.56 481.36 120.72 482.48 ;
      RECT 119.08 482.13 119.24 482.48 ;
      RECT 117.5 482.13 119.24 482.29 ;
      RECT 117.5 481.41 117.66 482.29 ;
      RECT 120.56 481.68 122.97 481.84 ;
      RECT 116.78 481.41 117.66 481.57 ;
      RECT 119.72 481.36 120.72 481.52 ;
      RECT 119.72 487.2 120.72 487.36 ;
      RECT 120.56 486.24 120.72 487.36 ;
      RECT 116.78 487.15 117.66 487.31 ;
      RECT 117.5 486.43 117.66 487.31 ;
      RECT 120.56 486.88 122.97 487.04 ;
      RECT 117.5 486.43 119.24 486.59 ;
      RECT 119.08 486.24 119.24 486.59 ;
      RECT 119.08 486.24 120.72 486.4 ;
      RECT 119.08 489.12 120.72 489.28 ;
      RECT 120.56 488.16 120.72 489.28 ;
      RECT 119.08 488.93 119.24 489.28 ;
      RECT 117.5 488.93 119.24 489.09 ;
      RECT 117.5 488.21 117.66 489.09 ;
      RECT 120.56 488.48 122.97 488.64 ;
      RECT 116.78 488.21 117.66 488.37 ;
      RECT 119.72 488.16 120.72 488.32 ;
      RECT 119.72 494 120.72 494.16 ;
      RECT 120.56 493.04 120.72 494.16 ;
      RECT 116.78 493.95 117.66 494.11 ;
      RECT 117.5 493.23 117.66 494.11 ;
      RECT 120.56 493.68 122.97 493.84 ;
      RECT 117.5 493.23 119.24 493.39 ;
      RECT 119.08 493.04 119.24 493.39 ;
      RECT 119.08 493.04 120.72 493.2 ;
      RECT 119.08 495.92 120.72 496.08 ;
      RECT 120.56 494.96 120.72 496.08 ;
      RECT 119.08 495.73 119.24 496.08 ;
      RECT 117.5 495.73 119.24 495.89 ;
      RECT 117.5 495.01 117.66 495.89 ;
      RECT 120.56 495.28 122.97 495.44 ;
      RECT 116.78 495.01 117.66 495.17 ;
      RECT 119.72 494.96 120.72 495.12 ;
      RECT 119.72 500.8 120.72 500.96 ;
      RECT 120.56 499.84 120.72 500.96 ;
      RECT 116.78 500.75 117.66 500.91 ;
      RECT 117.5 500.03 117.66 500.91 ;
      RECT 120.56 500.48 122.97 500.64 ;
      RECT 117.5 500.03 119.24 500.19 ;
      RECT 119.08 499.84 119.24 500.19 ;
      RECT 119.08 499.84 120.72 500 ;
      RECT 119.08 502.72 120.72 502.88 ;
      RECT 120.56 501.76 120.72 502.88 ;
      RECT 119.08 502.53 119.24 502.88 ;
      RECT 117.5 502.53 119.24 502.69 ;
      RECT 117.5 501.81 117.66 502.69 ;
      RECT 120.56 502.08 122.97 502.24 ;
      RECT 116.78 501.81 117.66 501.97 ;
      RECT 119.72 501.76 120.72 501.92 ;
      RECT 119.08 70.88 120.72 71.08 ;
      RECT 120.56 69.96 120.72 71.08 ;
      RECT 117.5 70.75 119.24 70.91 ;
      RECT 117.5 70.11 117.66 70.91 ;
      RECT 120.56 70.33 122.96 70.51 ;
      RECT 116.78 70.11 117.66 70.27 ;
      RECT 119.72 69.96 120.72 70.12 ;
      RECT 119.72 75.8 120.72 75.96 ;
      RECT 120.56 74.84 120.72 75.96 ;
      RECT 116.78 75.65 117.66 75.81 ;
      RECT 117.5 75.01 117.66 75.81 ;
      RECT 120.56 75.41 122.96 75.59 ;
      RECT 117.5 75.01 119.24 75.17 ;
      RECT 119.08 74.84 120.72 75.04 ;
      RECT 119.08 77.68 120.72 77.88 ;
      RECT 120.56 76.76 120.72 77.88 ;
      RECT 117.5 77.55 119.24 77.71 ;
      RECT 117.5 76.91 117.66 77.71 ;
      RECT 120.56 77.13 122.96 77.31 ;
      RECT 116.78 76.91 117.66 77.07 ;
      RECT 119.72 76.76 120.72 76.92 ;
      RECT 119.72 82.6 120.72 82.76 ;
      RECT 120.56 81.64 120.72 82.76 ;
      RECT 116.78 82.45 117.66 82.61 ;
      RECT 117.5 81.81 117.66 82.61 ;
      RECT 120.56 82.21 122.96 82.39 ;
      RECT 117.5 81.81 119.24 81.97 ;
      RECT 119.08 81.64 120.72 81.84 ;
      RECT 119.08 84.48 120.72 84.68 ;
      RECT 120.56 83.56 120.72 84.68 ;
      RECT 117.5 84.35 119.24 84.51 ;
      RECT 117.5 83.71 117.66 84.51 ;
      RECT 120.56 83.93 122.96 84.11 ;
      RECT 116.78 83.71 117.66 83.87 ;
      RECT 119.72 83.56 120.72 83.72 ;
      RECT 119.72 89.4 120.72 89.56 ;
      RECT 120.56 88.44 120.72 89.56 ;
      RECT 116.78 89.25 117.66 89.41 ;
      RECT 117.5 88.61 117.66 89.41 ;
      RECT 120.56 89.01 122.96 89.19 ;
      RECT 117.5 88.61 119.24 88.77 ;
      RECT 119.08 88.44 120.72 88.64 ;
      RECT 119.08 91.28 120.72 91.48 ;
      RECT 120.56 90.36 120.72 91.48 ;
      RECT 117.5 91.15 119.24 91.31 ;
      RECT 117.5 90.51 117.66 91.31 ;
      RECT 120.56 90.73 122.96 90.91 ;
      RECT 116.78 90.51 117.66 90.67 ;
      RECT 119.72 90.36 120.72 90.52 ;
      RECT 119.72 96.2 120.72 96.36 ;
      RECT 120.56 95.24 120.72 96.36 ;
      RECT 116.78 96.05 117.66 96.21 ;
      RECT 117.5 95.41 117.66 96.21 ;
      RECT 120.56 95.81 122.96 95.99 ;
      RECT 117.5 95.41 119.24 95.57 ;
      RECT 119.08 95.24 120.72 95.44 ;
      RECT 119.08 98.08 120.72 98.28 ;
      RECT 120.56 97.16 120.72 98.28 ;
      RECT 117.5 97.95 119.24 98.11 ;
      RECT 117.5 97.31 117.66 98.11 ;
      RECT 120.56 97.53 122.96 97.71 ;
      RECT 116.78 97.31 117.66 97.47 ;
      RECT 119.72 97.16 120.72 97.32 ;
      RECT 119.72 103 120.72 103.16 ;
      RECT 120.56 102.04 120.72 103.16 ;
      RECT 116.78 102.85 117.66 103.01 ;
      RECT 117.5 102.21 117.66 103.01 ;
      RECT 120.56 102.61 122.96 102.79 ;
      RECT 117.5 102.21 119.24 102.37 ;
      RECT 119.08 102.04 120.72 102.24 ;
      RECT 119.08 104.88 120.72 105.08 ;
      RECT 120.56 103.96 120.72 105.08 ;
      RECT 117.5 104.75 119.24 104.91 ;
      RECT 117.5 104.11 117.66 104.91 ;
      RECT 120.56 104.33 122.96 104.51 ;
      RECT 116.78 104.11 117.66 104.27 ;
      RECT 119.72 103.96 120.72 104.12 ;
      RECT 119.72 109.8 120.72 109.96 ;
      RECT 120.56 108.84 120.72 109.96 ;
      RECT 116.78 109.65 117.66 109.81 ;
      RECT 117.5 109.01 117.66 109.81 ;
      RECT 120.56 109.41 122.96 109.59 ;
      RECT 117.5 109.01 119.24 109.17 ;
      RECT 119.08 108.84 120.72 109.04 ;
      RECT 119.08 111.68 120.72 111.88 ;
      RECT 120.56 110.76 120.72 111.88 ;
      RECT 117.5 111.55 119.24 111.71 ;
      RECT 117.5 110.91 117.66 111.71 ;
      RECT 120.56 111.13 122.96 111.31 ;
      RECT 116.78 110.91 117.66 111.07 ;
      RECT 119.72 110.76 120.72 110.92 ;
      RECT 119.72 116.6 120.72 116.76 ;
      RECT 120.56 115.64 120.72 116.76 ;
      RECT 116.78 116.45 117.66 116.61 ;
      RECT 117.5 115.81 117.66 116.61 ;
      RECT 120.56 116.21 122.96 116.39 ;
      RECT 117.5 115.81 119.24 115.97 ;
      RECT 119.08 115.64 120.72 115.84 ;
      RECT 119.08 118.48 120.72 118.68 ;
      RECT 120.56 117.56 120.72 118.68 ;
      RECT 117.5 118.35 119.24 118.51 ;
      RECT 117.5 117.71 117.66 118.51 ;
      RECT 120.56 117.93 122.96 118.11 ;
      RECT 116.78 117.71 117.66 117.87 ;
      RECT 119.72 117.56 120.72 117.72 ;
      RECT 119.72 123.4 120.72 123.56 ;
      RECT 120.56 122.44 120.72 123.56 ;
      RECT 116.78 123.25 117.66 123.41 ;
      RECT 117.5 122.61 117.66 123.41 ;
      RECT 120.56 123.01 122.96 123.19 ;
      RECT 117.5 122.61 119.24 122.77 ;
      RECT 119.08 122.44 120.72 122.64 ;
      RECT 119.08 125.28 120.72 125.48 ;
      RECT 120.56 124.36 120.72 125.48 ;
      RECT 117.5 125.15 119.24 125.31 ;
      RECT 117.5 124.51 117.66 125.31 ;
      RECT 120.56 124.73 122.96 124.91 ;
      RECT 116.78 124.51 117.66 124.67 ;
      RECT 119.72 124.36 120.72 124.52 ;
      RECT 119.72 130.2 120.72 130.36 ;
      RECT 120.56 129.24 120.72 130.36 ;
      RECT 116.78 130.05 117.66 130.21 ;
      RECT 117.5 129.41 117.66 130.21 ;
      RECT 120.56 129.81 122.96 129.99 ;
      RECT 117.5 129.41 119.24 129.57 ;
      RECT 119.08 129.24 120.72 129.44 ;
      RECT 119.08 132.08 120.72 132.28 ;
      RECT 120.56 131.16 120.72 132.28 ;
      RECT 117.5 131.95 119.24 132.11 ;
      RECT 117.5 131.31 117.66 132.11 ;
      RECT 120.56 131.53 122.96 131.71 ;
      RECT 116.78 131.31 117.66 131.47 ;
      RECT 119.72 131.16 120.72 131.32 ;
      RECT 119.72 137 120.72 137.16 ;
      RECT 120.56 136.04 120.72 137.16 ;
      RECT 116.78 136.85 117.66 137.01 ;
      RECT 117.5 136.21 117.66 137.01 ;
      RECT 120.56 136.61 122.96 136.79 ;
      RECT 117.5 136.21 119.24 136.37 ;
      RECT 119.08 136.04 120.72 136.24 ;
      RECT 119.08 138.88 120.72 139.08 ;
      RECT 120.56 137.96 120.72 139.08 ;
      RECT 117.5 138.75 119.24 138.91 ;
      RECT 117.5 138.11 117.66 138.91 ;
      RECT 120.56 138.33 122.96 138.51 ;
      RECT 116.78 138.11 117.66 138.27 ;
      RECT 119.72 137.96 120.72 138.12 ;
      RECT 119.72 143.8 120.72 143.96 ;
      RECT 120.56 142.84 120.72 143.96 ;
      RECT 116.78 143.65 117.66 143.81 ;
      RECT 117.5 143.01 117.66 143.81 ;
      RECT 120.56 143.41 122.96 143.59 ;
      RECT 117.5 143.01 119.24 143.17 ;
      RECT 119.08 142.84 120.72 143.04 ;
      RECT 119.08 145.68 120.72 145.88 ;
      RECT 120.56 144.76 120.72 145.88 ;
      RECT 117.5 145.55 119.24 145.71 ;
      RECT 117.5 144.91 117.66 145.71 ;
      RECT 120.56 145.13 122.96 145.31 ;
      RECT 116.78 144.91 117.66 145.07 ;
      RECT 119.72 144.76 120.72 144.92 ;
      RECT 119.72 150.6 120.72 150.76 ;
      RECT 120.56 149.64 120.72 150.76 ;
      RECT 116.78 150.45 117.66 150.61 ;
      RECT 117.5 149.81 117.66 150.61 ;
      RECT 120.56 150.21 122.96 150.39 ;
      RECT 117.5 149.81 119.24 149.97 ;
      RECT 119.08 149.64 120.72 149.84 ;
      RECT 119.08 152.48 120.72 152.68 ;
      RECT 120.56 151.56 120.72 152.68 ;
      RECT 117.5 152.35 119.24 152.51 ;
      RECT 117.5 151.71 117.66 152.51 ;
      RECT 120.56 151.93 122.96 152.11 ;
      RECT 116.78 151.71 117.66 151.87 ;
      RECT 119.72 151.56 120.72 151.72 ;
      RECT 119.72 157.4 120.72 157.56 ;
      RECT 120.56 156.44 120.72 157.56 ;
      RECT 116.78 157.25 117.66 157.41 ;
      RECT 117.5 156.61 117.66 157.41 ;
      RECT 120.56 157.01 122.96 157.19 ;
      RECT 117.5 156.61 119.24 156.77 ;
      RECT 119.08 156.44 120.72 156.64 ;
      RECT 119.08 159.28 120.72 159.48 ;
      RECT 120.56 158.36 120.72 159.48 ;
      RECT 117.5 159.15 119.24 159.31 ;
      RECT 117.5 158.51 117.66 159.31 ;
      RECT 120.56 158.73 122.96 158.91 ;
      RECT 116.78 158.51 117.66 158.67 ;
      RECT 119.72 158.36 120.72 158.52 ;
      RECT 119.72 164.2 120.72 164.36 ;
      RECT 120.56 163.24 120.72 164.36 ;
      RECT 116.78 164.05 117.66 164.21 ;
      RECT 117.5 163.41 117.66 164.21 ;
      RECT 120.56 163.81 122.96 163.99 ;
      RECT 117.5 163.41 119.24 163.57 ;
      RECT 119.08 163.24 120.72 163.44 ;
      RECT 119.08 166.08 120.72 166.28 ;
      RECT 120.56 165.16 120.72 166.28 ;
      RECT 117.5 165.95 119.24 166.11 ;
      RECT 117.5 165.31 117.66 166.11 ;
      RECT 120.56 165.53 122.96 165.71 ;
      RECT 116.78 165.31 117.66 165.47 ;
      RECT 119.72 165.16 120.72 165.32 ;
      RECT 119.72 171 120.72 171.16 ;
      RECT 120.56 170.04 120.72 171.16 ;
      RECT 116.78 170.85 117.66 171.01 ;
      RECT 117.5 170.21 117.66 171.01 ;
      RECT 120.56 170.61 122.96 170.79 ;
      RECT 117.5 170.21 119.24 170.37 ;
      RECT 119.08 170.04 120.72 170.24 ;
      RECT 119.08 172.88 120.72 173.08 ;
      RECT 120.56 171.96 120.72 173.08 ;
      RECT 117.5 172.75 119.24 172.91 ;
      RECT 117.5 172.11 117.66 172.91 ;
      RECT 120.56 172.33 122.96 172.51 ;
      RECT 116.78 172.11 117.66 172.27 ;
      RECT 119.72 171.96 120.72 172.12 ;
      RECT 119.72 177.8 120.72 177.96 ;
      RECT 120.56 176.84 120.72 177.96 ;
      RECT 116.78 177.65 117.66 177.81 ;
      RECT 117.5 177.01 117.66 177.81 ;
      RECT 120.56 177.41 122.96 177.59 ;
      RECT 117.5 177.01 119.24 177.17 ;
      RECT 119.08 176.84 120.72 177.04 ;
      RECT 119.08 179.68 120.72 179.88 ;
      RECT 120.56 178.76 120.72 179.88 ;
      RECT 117.5 179.55 119.24 179.71 ;
      RECT 117.5 178.91 117.66 179.71 ;
      RECT 120.56 179.13 122.96 179.31 ;
      RECT 116.78 178.91 117.66 179.07 ;
      RECT 119.72 178.76 120.72 178.92 ;
      RECT 119.72 184.6 120.72 184.76 ;
      RECT 120.56 183.64 120.72 184.76 ;
      RECT 116.78 184.45 117.66 184.61 ;
      RECT 117.5 183.81 117.66 184.61 ;
      RECT 120.56 184.21 122.96 184.39 ;
      RECT 117.5 183.81 119.24 183.97 ;
      RECT 119.08 183.64 120.72 183.84 ;
      RECT 119.08 186.48 120.72 186.68 ;
      RECT 120.56 185.56 120.72 186.68 ;
      RECT 117.5 186.35 119.24 186.51 ;
      RECT 117.5 185.71 117.66 186.51 ;
      RECT 120.56 185.93 122.96 186.11 ;
      RECT 116.78 185.71 117.66 185.87 ;
      RECT 119.72 185.56 120.72 185.72 ;
      RECT 119.72 191.4 120.72 191.56 ;
      RECT 120.56 190.44 120.72 191.56 ;
      RECT 116.78 191.25 117.66 191.41 ;
      RECT 117.5 190.61 117.66 191.41 ;
      RECT 120.56 191.01 122.96 191.19 ;
      RECT 117.5 190.61 119.24 190.77 ;
      RECT 119.08 190.44 120.72 190.64 ;
      RECT 119.08 193.28 120.72 193.48 ;
      RECT 120.56 192.36 120.72 193.48 ;
      RECT 117.5 193.15 119.24 193.31 ;
      RECT 117.5 192.51 117.66 193.31 ;
      RECT 120.56 192.73 122.96 192.91 ;
      RECT 116.78 192.51 117.66 192.67 ;
      RECT 119.72 192.36 120.72 192.52 ;
      RECT 119.72 198.2 120.72 198.36 ;
      RECT 120.56 197.24 120.72 198.36 ;
      RECT 116.78 198.05 117.66 198.21 ;
      RECT 117.5 197.41 117.66 198.21 ;
      RECT 120.56 197.81 122.96 197.99 ;
      RECT 117.5 197.41 119.24 197.57 ;
      RECT 119.08 197.24 120.72 197.44 ;
      RECT 119.08 200.08 120.72 200.28 ;
      RECT 120.56 199.16 120.72 200.28 ;
      RECT 117.5 199.95 119.24 200.11 ;
      RECT 117.5 199.31 117.66 200.11 ;
      RECT 120.56 199.53 122.96 199.71 ;
      RECT 116.78 199.31 117.66 199.47 ;
      RECT 119.72 199.16 120.72 199.32 ;
      RECT 119.72 205 120.72 205.16 ;
      RECT 120.56 204.04 120.72 205.16 ;
      RECT 116.78 204.85 117.66 205.01 ;
      RECT 117.5 204.21 117.66 205.01 ;
      RECT 120.56 204.61 122.96 204.79 ;
      RECT 117.5 204.21 119.24 204.37 ;
      RECT 119.08 204.04 120.72 204.24 ;
      RECT 119.08 206.88 120.72 207.08 ;
      RECT 120.56 205.96 120.72 207.08 ;
      RECT 117.5 206.75 119.24 206.91 ;
      RECT 117.5 206.11 117.66 206.91 ;
      RECT 120.56 206.33 122.96 206.51 ;
      RECT 116.78 206.11 117.66 206.27 ;
      RECT 119.72 205.96 120.72 206.12 ;
      RECT 119.72 211.8 120.72 211.96 ;
      RECT 120.56 210.84 120.72 211.96 ;
      RECT 116.78 211.65 117.66 211.81 ;
      RECT 117.5 211.01 117.66 211.81 ;
      RECT 120.56 211.41 122.96 211.59 ;
      RECT 117.5 211.01 119.24 211.17 ;
      RECT 119.08 210.84 120.72 211.04 ;
      RECT 119.08 213.68 120.72 213.88 ;
      RECT 120.56 212.76 120.72 213.88 ;
      RECT 117.5 213.55 119.24 213.71 ;
      RECT 117.5 212.91 117.66 213.71 ;
      RECT 120.56 213.13 122.96 213.31 ;
      RECT 116.78 212.91 117.66 213.07 ;
      RECT 119.72 212.76 120.72 212.92 ;
      RECT 119.72 218.6 120.72 218.76 ;
      RECT 120.56 217.64 120.72 218.76 ;
      RECT 116.78 218.45 117.66 218.61 ;
      RECT 117.5 217.81 117.66 218.61 ;
      RECT 120.56 218.21 122.96 218.39 ;
      RECT 117.5 217.81 119.24 217.97 ;
      RECT 119.08 217.64 120.72 217.84 ;
      RECT 119.08 220.48 120.72 220.68 ;
      RECT 120.56 219.56 120.72 220.68 ;
      RECT 117.5 220.35 119.24 220.51 ;
      RECT 117.5 219.71 117.66 220.51 ;
      RECT 120.56 219.93 122.96 220.11 ;
      RECT 116.78 219.71 117.66 219.87 ;
      RECT 119.72 219.56 120.72 219.72 ;
      RECT 119.72 225.4 120.72 225.56 ;
      RECT 120.56 224.44 120.72 225.56 ;
      RECT 116.78 225.25 117.66 225.41 ;
      RECT 117.5 224.61 117.66 225.41 ;
      RECT 120.56 225.01 122.96 225.19 ;
      RECT 117.5 224.61 119.24 224.77 ;
      RECT 119.08 224.44 120.72 224.64 ;
      RECT 119.08 227.28 120.72 227.48 ;
      RECT 120.56 226.36 120.72 227.48 ;
      RECT 117.5 227.15 119.24 227.31 ;
      RECT 117.5 226.51 117.66 227.31 ;
      RECT 120.56 226.73 122.96 226.91 ;
      RECT 116.78 226.51 117.66 226.67 ;
      RECT 119.72 226.36 120.72 226.52 ;
      RECT 119.72 232.2 120.72 232.36 ;
      RECT 120.56 231.24 120.72 232.36 ;
      RECT 116.78 232.05 117.66 232.21 ;
      RECT 117.5 231.41 117.66 232.21 ;
      RECT 120.56 231.81 122.96 231.99 ;
      RECT 117.5 231.41 119.24 231.57 ;
      RECT 119.08 231.24 120.72 231.44 ;
      RECT 119.08 234.08 120.72 234.28 ;
      RECT 120.56 233.16 120.72 234.28 ;
      RECT 117.5 233.95 119.24 234.11 ;
      RECT 117.5 233.31 117.66 234.11 ;
      RECT 120.56 233.53 122.96 233.71 ;
      RECT 116.78 233.31 117.66 233.47 ;
      RECT 119.72 233.16 120.72 233.32 ;
      RECT 119.72 239 120.72 239.16 ;
      RECT 120.56 238.04 120.72 239.16 ;
      RECT 116.78 238.85 117.66 239.01 ;
      RECT 117.5 238.21 117.66 239.01 ;
      RECT 120.56 238.61 122.96 238.79 ;
      RECT 117.5 238.21 119.24 238.37 ;
      RECT 119.08 238.04 120.72 238.24 ;
      RECT 119.08 240.88 120.72 241.08 ;
      RECT 120.56 239.96 120.72 241.08 ;
      RECT 117.5 240.75 119.24 240.91 ;
      RECT 117.5 240.11 117.66 240.91 ;
      RECT 120.56 240.33 122.96 240.51 ;
      RECT 116.78 240.11 117.66 240.27 ;
      RECT 119.72 239.96 120.72 240.12 ;
      RECT 119.72 245.8 120.72 245.96 ;
      RECT 120.56 244.84 120.72 245.96 ;
      RECT 116.78 245.65 117.66 245.81 ;
      RECT 117.5 245.01 117.66 245.81 ;
      RECT 120.56 245.41 122.96 245.59 ;
      RECT 117.5 245.01 119.24 245.17 ;
      RECT 119.08 244.84 120.72 245.04 ;
      RECT 119.08 247.68 120.72 247.88 ;
      RECT 120.56 246.76 120.72 247.88 ;
      RECT 117.5 247.55 119.24 247.71 ;
      RECT 117.5 246.91 117.66 247.71 ;
      RECT 120.56 247.13 122.96 247.31 ;
      RECT 116.78 246.91 117.66 247.07 ;
      RECT 119.72 246.76 120.72 246.92 ;
      RECT 119.72 252.6 120.72 252.76 ;
      RECT 120.56 251.64 120.72 252.76 ;
      RECT 116.78 252.45 117.66 252.61 ;
      RECT 117.5 251.81 117.66 252.61 ;
      RECT 120.56 252.21 122.96 252.39 ;
      RECT 117.5 251.81 119.24 251.97 ;
      RECT 119.08 251.64 120.72 251.84 ;
      RECT 119.08 254.48 120.72 254.68 ;
      RECT 120.56 253.56 120.72 254.68 ;
      RECT 117.5 254.35 119.24 254.51 ;
      RECT 117.5 253.71 117.66 254.51 ;
      RECT 120.56 253.93 122.96 254.11 ;
      RECT 116.78 253.71 117.66 253.87 ;
      RECT 119.72 253.56 120.72 253.72 ;
      RECT 119.72 259.4 120.72 259.56 ;
      RECT 120.56 258.44 120.72 259.56 ;
      RECT 116.78 259.25 117.66 259.41 ;
      RECT 117.5 258.61 117.66 259.41 ;
      RECT 120.56 259.01 122.96 259.19 ;
      RECT 117.5 258.61 119.24 258.77 ;
      RECT 119.08 258.44 120.72 258.64 ;
      RECT 119.08 261.28 120.72 261.48 ;
      RECT 120.56 260.36 120.72 261.48 ;
      RECT 117.5 261.15 119.24 261.31 ;
      RECT 117.5 260.51 117.66 261.31 ;
      RECT 120.56 260.73 122.96 260.91 ;
      RECT 116.78 260.51 117.66 260.67 ;
      RECT 119.72 260.36 120.72 260.52 ;
      RECT 119.72 266.2 120.72 266.36 ;
      RECT 120.56 265.24 120.72 266.36 ;
      RECT 116.78 266.05 117.66 266.21 ;
      RECT 117.5 265.41 117.66 266.21 ;
      RECT 120.56 265.81 122.96 265.99 ;
      RECT 117.5 265.41 119.24 265.57 ;
      RECT 119.08 265.24 120.72 265.44 ;
      RECT 119.08 268.08 120.72 268.28 ;
      RECT 120.56 267.16 120.72 268.28 ;
      RECT 117.5 267.95 119.24 268.11 ;
      RECT 117.5 267.31 117.66 268.11 ;
      RECT 120.56 267.53 122.96 267.71 ;
      RECT 116.78 267.31 117.66 267.47 ;
      RECT 119.72 267.16 120.72 267.32 ;
      RECT 119.72 273 120.72 273.16 ;
      RECT 120.56 272.04 120.72 273.16 ;
      RECT 116.78 272.85 117.66 273.01 ;
      RECT 117.5 272.21 117.66 273.01 ;
      RECT 120.56 272.61 122.96 272.79 ;
      RECT 117.5 272.21 119.24 272.37 ;
      RECT 119.08 272.04 120.72 272.24 ;
      RECT 119.08 274.88 120.72 275.08 ;
      RECT 120.56 273.96 120.72 275.08 ;
      RECT 117.5 274.75 119.24 274.91 ;
      RECT 117.5 274.11 117.66 274.91 ;
      RECT 120.56 274.33 122.96 274.51 ;
      RECT 116.78 274.11 117.66 274.27 ;
      RECT 119.72 273.96 120.72 274.12 ;
      RECT 119.72 279.8 120.72 279.96 ;
      RECT 120.56 278.84 120.72 279.96 ;
      RECT 116.78 279.65 117.66 279.81 ;
      RECT 117.5 279.01 117.66 279.81 ;
      RECT 120.56 279.41 122.96 279.59 ;
      RECT 117.5 279.01 119.24 279.17 ;
      RECT 119.08 278.84 120.72 279.04 ;
      RECT 119.08 281.68 120.72 281.88 ;
      RECT 120.56 280.76 120.72 281.88 ;
      RECT 117.5 281.55 119.24 281.71 ;
      RECT 117.5 280.91 117.66 281.71 ;
      RECT 120.56 281.13 122.96 281.31 ;
      RECT 116.78 280.91 117.66 281.07 ;
      RECT 119.72 280.76 120.72 280.92 ;
      RECT 119.72 286.6 120.72 286.76 ;
      RECT 120.56 285.64 120.72 286.76 ;
      RECT 116.78 286.45 117.66 286.61 ;
      RECT 117.5 285.81 117.66 286.61 ;
      RECT 120.56 286.21 122.96 286.39 ;
      RECT 117.5 285.81 119.24 285.97 ;
      RECT 119.08 285.64 120.72 285.84 ;
      RECT 119.08 288.48 120.72 288.68 ;
      RECT 120.56 287.56 120.72 288.68 ;
      RECT 117.5 288.35 119.24 288.51 ;
      RECT 117.5 287.71 117.66 288.51 ;
      RECT 120.56 287.93 122.96 288.11 ;
      RECT 116.78 287.71 117.66 287.87 ;
      RECT 119.72 287.56 120.72 287.72 ;
      RECT 119.72 293.4 120.72 293.56 ;
      RECT 120.56 292.44 120.72 293.56 ;
      RECT 116.78 293.25 117.66 293.41 ;
      RECT 117.5 292.61 117.66 293.41 ;
      RECT 120.56 293.01 122.96 293.19 ;
      RECT 117.5 292.61 119.24 292.77 ;
      RECT 119.08 292.44 120.72 292.64 ;
      RECT 119.08 295.28 120.72 295.48 ;
      RECT 120.56 294.36 120.72 295.48 ;
      RECT 117.5 295.15 119.24 295.31 ;
      RECT 117.5 294.51 117.66 295.31 ;
      RECT 120.56 294.73 122.96 294.91 ;
      RECT 116.78 294.51 117.66 294.67 ;
      RECT 119.72 294.36 120.72 294.52 ;
      RECT 119.72 300.2 120.72 300.36 ;
      RECT 120.56 299.24 120.72 300.36 ;
      RECT 116.78 300.05 117.66 300.21 ;
      RECT 117.5 299.41 117.66 300.21 ;
      RECT 120.56 299.81 122.96 299.99 ;
      RECT 117.5 299.41 119.24 299.57 ;
      RECT 119.08 299.24 120.72 299.44 ;
      RECT 119.08 302.08 120.72 302.28 ;
      RECT 120.56 301.16 120.72 302.28 ;
      RECT 117.5 301.95 119.24 302.11 ;
      RECT 117.5 301.31 117.66 302.11 ;
      RECT 120.56 301.53 122.96 301.71 ;
      RECT 116.78 301.31 117.66 301.47 ;
      RECT 119.72 301.16 120.72 301.32 ;
      RECT 119.72 307 120.72 307.16 ;
      RECT 120.56 306.04 120.72 307.16 ;
      RECT 116.78 306.85 117.66 307.01 ;
      RECT 117.5 306.21 117.66 307.01 ;
      RECT 120.56 306.61 122.96 306.79 ;
      RECT 117.5 306.21 119.24 306.37 ;
      RECT 119.08 306.04 120.72 306.24 ;
      RECT 119.08 308.88 120.72 309.08 ;
      RECT 120.56 307.96 120.72 309.08 ;
      RECT 117.5 308.75 119.24 308.91 ;
      RECT 117.5 308.11 117.66 308.91 ;
      RECT 120.56 308.33 122.96 308.51 ;
      RECT 116.78 308.11 117.66 308.27 ;
      RECT 119.72 307.96 120.72 308.12 ;
      RECT 119.72 313.8 120.72 313.96 ;
      RECT 120.56 312.84 120.72 313.96 ;
      RECT 116.78 313.65 117.66 313.81 ;
      RECT 117.5 313.01 117.66 313.81 ;
      RECT 120.56 313.41 122.96 313.59 ;
      RECT 117.5 313.01 119.24 313.17 ;
      RECT 119.08 312.84 120.72 313.04 ;
      RECT 119.08 315.68 120.72 315.88 ;
      RECT 120.56 314.76 120.72 315.88 ;
      RECT 117.5 315.55 119.24 315.71 ;
      RECT 117.5 314.91 117.66 315.71 ;
      RECT 120.56 315.13 122.96 315.31 ;
      RECT 116.78 314.91 117.66 315.07 ;
      RECT 119.72 314.76 120.72 314.92 ;
      RECT 119.72 320.6 120.72 320.76 ;
      RECT 120.56 319.64 120.72 320.76 ;
      RECT 116.78 320.45 117.66 320.61 ;
      RECT 117.5 319.81 117.66 320.61 ;
      RECT 120.56 320.21 122.96 320.39 ;
      RECT 117.5 319.81 119.24 319.97 ;
      RECT 119.08 319.64 120.72 319.84 ;
      RECT 119.08 322.48 120.72 322.68 ;
      RECT 120.56 321.56 120.72 322.68 ;
      RECT 117.5 322.35 119.24 322.51 ;
      RECT 117.5 321.71 117.66 322.51 ;
      RECT 120.56 321.93 122.96 322.11 ;
      RECT 116.78 321.71 117.66 321.87 ;
      RECT 119.72 321.56 120.72 321.72 ;
      RECT 119.72 327.4 120.72 327.56 ;
      RECT 120.56 326.44 120.72 327.56 ;
      RECT 116.78 327.25 117.66 327.41 ;
      RECT 117.5 326.61 117.66 327.41 ;
      RECT 120.56 327.01 122.96 327.19 ;
      RECT 117.5 326.61 119.24 326.77 ;
      RECT 119.08 326.44 120.72 326.64 ;
      RECT 119.08 329.28 120.72 329.48 ;
      RECT 120.56 328.36 120.72 329.48 ;
      RECT 117.5 329.15 119.24 329.31 ;
      RECT 117.5 328.51 117.66 329.31 ;
      RECT 120.56 328.73 122.96 328.91 ;
      RECT 116.78 328.51 117.66 328.67 ;
      RECT 119.72 328.36 120.72 328.52 ;
      RECT 119.72 334.2 120.72 334.36 ;
      RECT 120.56 333.24 120.72 334.36 ;
      RECT 116.78 334.05 117.66 334.21 ;
      RECT 117.5 333.41 117.66 334.21 ;
      RECT 120.56 333.81 122.96 333.99 ;
      RECT 117.5 333.41 119.24 333.57 ;
      RECT 119.08 333.24 120.72 333.44 ;
      RECT 119.08 336.08 120.72 336.28 ;
      RECT 120.56 335.16 120.72 336.28 ;
      RECT 117.5 335.95 119.24 336.11 ;
      RECT 117.5 335.31 117.66 336.11 ;
      RECT 120.56 335.53 122.96 335.71 ;
      RECT 116.78 335.31 117.66 335.47 ;
      RECT 119.72 335.16 120.72 335.32 ;
      RECT 119.72 341 120.72 341.16 ;
      RECT 120.56 340.04 120.72 341.16 ;
      RECT 116.78 340.85 117.66 341.01 ;
      RECT 117.5 340.21 117.66 341.01 ;
      RECT 120.56 340.61 122.96 340.79 ;
      RECT 117.5 340.21 119.24 340.37 ;
      RECT 119.08 340.04 120.72 340.24 ;
      RECT 119.08 342.88 120.72 343.08 ;
      RECT 120.56 341.96 120.72 343.08 ;
      RECT 117.5 342.75 119.24 342.91 ;
      RECT 117.5 342.11 117.66 342.91 ;
      RECT 120.56 342.33 122.96 342.51 ;
      RECT 116.78 342.11 117.66 342.27 ;
      RECT 119.72 341.96 120.72 342.12 ;
      RECT 119.72 347.8 120.72 347.96 ;
      RECT 120.56 346.84 120.72 347.96 ;
      RECT 116.78 347.65 117.66 347.81 ;
      RECT 117.5 347.01 117.66 347.81 ;
      RECT 120.56 347.41 122.96 347.59 ;
      RECT 117.5 347.01 119.24 347.17 ;
      RECT 119.08 346.84 120.72 347.04 ;
      RECT 119.08 349.68 120.72 349.88 ;
      RECT 120.56 348.76 120.72 349.88 ;
      RECT 117.5 349.55 119.24 349.71 ;
      RECT 117.5 348.91 117.66 349.71 ;
      RECT 120.56 349.13 122.96 349.31 ;
      RECT 116.78 348.91 117.66 349.07 ;
      RECT 119.72 348.76 120.72 348.92 ;
      RECT 119.72 354.6 120.72 354.76 ;
      RECT 120.56 353.64 120.72 354.76 ;
      RECT 116.78 354.45 117.66 354.61 ;
      RECT 117.5 353.81 117.66 354.61 ;
      RECT 120.56 354.21 122.96 354.39 ;
      RECT 117.5 353.81 119.24 353.97 ;
      RECT 119.08 353.64 120.72 353.84 ;
      RECT 119.08 356.48 120.72 356.68 ;
      RECT 120.56 355.56 120.72 356.68 ;
      RECT 117.5 356.35 119.24 356.51 ;
      RECT 117.5 355.71 117.66 356.51 ;
      RECT 120.56 355.93 122.96 356.11 ;
      RECT 116.78 355.71 117.66 355.87 ;
      RECT 119.72 355.56 120.72 355.72 ;
      RECT 119.72 361.4 120.72 361.56 ;
      RECT 120.56 360.44 120.72 361.56 ;
      RECT 116.78 361.25 117.66 361.41 ;
      RECT 117.5 360.61 117.66 361.41 ;
      RECT 120.56 361.01 122.96 361.19 ;
      RECT 117.5 360.61 119.24 360.77 ;
      RECT 119.08 360.44 120.72 360.64 ;
      RECT 119.08 363.28 120.72 363.48 ;
      RECT 120.56 362.36 120.72 363.48 ;
      RECT 117.5 363.15 119.24 363.31 ;
      RECT 117.5 362.51 117.66 363.31 ;
      RECT 120.56 362.73 122.96 362.91 ;
      RECT 116.78 362.51 117.66 362.67 ;
      RECT 119.72 362.36 120.72 362.52 ;
      RECT 119.72 368.2 120.72 368.36 ;
      RECT 120.56 367.24 120.72 368.36 ;
      RECT 116.78 368.05 117.66 368.21 ;
      RECT 117.5 367.41 117.66 368.21 ;
      RECT 120.56 367.81 122.96 367.99 ;
      RECT 117.5 367.41 119.24 367.57 ;
      RECT 119.08 367.24 120.72 367.44 ;
      RECT 119.08 370.08 120.72 370.28 ;
      RECT 120.56 369.16 120.72 370.28 ;
      RECT 117.5 369.95 119.24 370.11 ;
      RECT 117.5 369.31 117.66 370.11 ;
      RECT 120.56 369.53 122.96 369.71 ;
      RECT 116.78 369.31 117.66 369.47 ;
      RECT 119.72 369.16 120.72 369.32 ;
      RECT 119.72 375 120.72 375.16 ;
      RECT 120.56 374.04 120.72 375.16 ;
      RECT 116.78 374.85 117.66 375.01 ;
      RECT 117.5 374.21 117.66 375.01 ;
      RECT 120.56 374.61 122.96 374.79 ;
      RECT 117.5 374.21 119.24 374.37 ;
      RECT 119.08 374.04 120.72 374.24 ;
      RECT 119.08 376.88 120.72 377.08 ;
      RECT 120.56 375.96 120.72 377.08 ;
      RECT 117.5 376.75 119.24 376.91 ;
      RECT 117.5 376.11 117.66 376.91 ;
      RECT 120.56 376.33 122.96 376.51 ;
      RECT 116.78 376.11 117.66 376.27 ;
      RECT 119.72 375.96 120.72 376.12 ;
      RECT 119.72 381.8 120.72 381.96 ;
      RECT 120.56 380.84 120.72 381.96 ;
      RECT 116.78 381.65 117.66 381.81 ;
      RECT 117.5 381.01 117.66 381.81 ;
      RECT 120.56 381.41 122.96 381.59 ;
      RECT 117.5 381.01 119.24 381.17 ;
      RECT 119.08 380.84 120.72 381.04 ;
      RECT 119.08 383.68 120.72 383.88 ;
      RECT 120.56 382.76 120.72 383.88 ;
      RECT 117.5 383.55 119.24 383.71 ;
      RECT 117.5 382.91 117.66 383.71 ;
      RECT 120.56 383.13 122.96 383.31 ;
      RECT 116.78 382.91 117.66 383.07 ;
      RECT 119.72 382.76 120.72 382.92 ;
      RECT 119.72 388.6 120.72 388.76 ;
      RECT 120.56 387.64 120.72 388.76 ;
      RECT 116.78 388.45 117.66 388.61 ;
      RECT 117.5 387.81 117.66 388.61 ;
      RECT 120.56 388.21 122.96 388.39 ;
      RECT 117.5 387.81 119.24 387.97 ;
      RECT 119.08 387.64 120.72 387.84 ;
      RECT 119.08 390.48 120.72 390.68 ;
      RECT 120.56 389.56 120.72 390.68 ;
      RECT 117.5 390.35 119.24 390.51 ;
      RECT 117.5 389.71 117.66 390.51 ;
      RECT 120.56 389.93 122.96 390.11 ;
      RECT 116.78 389.71 117.66 389.87 ;
      RECT 119.72 389.56 120.72 389.72 ;
      RECT 119.72 395.4 120.72 395.56 ;
      RECT 120.56 394.44 120.72 395.56 ;
      RECT 116.78 395.25 117.66 395.41 ;
      RECT 117.5 394.61 117.66 395.41 ;
      RECT 120.56 395.01 122.96 395.19 ;
      RECT 117.5 394.61 119.24 394.77 ;
      RECT 119.08 394.44 120.72 394.64 ;
      RECT 119.08 397.28 120.72 397.48 ;
      RECT 120.56 396.36 120.72 397.48 ;
      RECT 117.5 397.15 119.24 397.31 ;
      RECT 117.5 396.51 117.66 397.31 ;
      RECT 120.56 396.73 122.96 396.91 ;
      RECT 116.78 396.51 117.66 396.67 ;
      RECT 119.72 396.36 120.72 396.52 ;
      RECT 119.72 402.2 120.72 402.36 ;
      RECT 120.56 401.24 120.72 402.36 ;
      RECT 116.78 402.05 117.66 402.21 ;
      RECT 117.5 401.41 117.66 402.21 ;
      RECT 120.56 401.81 122.96 401.99 ;
      RECT 117.5 401.41 119.24 401.57 ;
      RECT 119.08 401.24 120.72 401.44 ;
      RECT 119.08 404.08 120.72 404.28 ;
      RECT 120.56 403.16 120.72 404.28 ;
      RECT 117.5 403.95 119.24 404.11 ;
      RECT 117.5 403.31 117.66 404.11 ;
      RECT 120.56 403.53 122.96 403.71 ;
      RECT 116.78 403.31 117.66 403.47 ;
      RECT 119.72 403.16 120.72 403.32 ;
      RECT 119.72 409 120.72 409.16 ;
      RECT 120.56 408.04 120.72 409.16 ;
      RECT 116.78 408.85 117.66 409.01 ;
      RECT 117.5 408.21 117.66 409.01 ;
      RECT 120.56 408.61 122.96 408.79 ;
      RECT 117.5 408.21 119.24 408.37 ;
      RECT 119.08 408.04 120.72 408.24 ;
      RECT 119.08 410.88 120.72 411.08 ;
      RECT 120.56 409.96 120.72 411.08 ;
      RECT 117.5 410.75 119.24 410.91 ;
      RECT 117.5 410.11 117.66 410.91 ;
      RECT 120.56 410.33 122.96 410.51 ;
      RECT 116.78 410.11 117.66 410.27 ;
      RECT 119.72 409.96 120.72 410.12 ;
      RECT 119.72 415.8 120.72 415.96 ;
      RECT 120.56 414.84 120.72 415.96 ;
      RECT 116.78 415.65 117.66 415.81 ;
      RECT 117.5 415.01 117.66 415.81 ;
      RECT 120.56 415.41 122.96 415.59 ;
      RECT 117.5 415.01 119.24 415.17 ;
      RECT 119.08 414.84 120.72 415.04 ;
      RECT 119.08 417.68 120.72 417.88 ;
      RECT 120.56 416.76 120.72 417.88 ;
      RECT 117.5 417.55 119.24 417.71 ;
      RECT 117.5 416.91 117.66 417.71 ;
      RECT 120.56 417.13 122.96 417.31 ;
      RECT 116.78 416.91 117.66 417.07 ;
      RECT 119.72 416.76 120.72 416.92 ;
      RECT 119.72 422.6 120.72 422.76 ;
      RECT 120.56 421.64 120.72 422.76 ;
      RECT 116.78 422.45 117.66 422.61 ;
      RECT 117.5 421.81 117.66 422.61 ;
      RECT 120.56 422.21 122.96 422.39 ;
      RECT 117.5 421.81 119.24 421.97 ;
      RECT 119.08 421.64 120.72 421.84 ;
      RECT 119.08 424.48 120.72 424.68 ;
      RECT 120.56 423.56 120.72 424.68 ;
      RECT 117.5 424.35 119.24 424.51 ;
      RECT 117.5 423.71 117.66 424.51 ;
      RECT 120.56 423.93 122.96 424.11 ;
      RECT 116.78 423.71 117.66 423.87 ;
      RECT 119.72 423.56 120.72 423.72 ;
      RECT 119.72 429.4 120.72 429.56 ;
      RECT 120.56 428.44 120.72 429.56 ;
      RECT 116.78 429.25 117.66 429.41 ;
      RECT 117.5 428.61 117.66 429.41 ;
      RECT 120.56 429.01 122.96 429.19 ;
      RECT 117.5 428.61 119.24 428.77 ;
      RECT 119.08 428.44 120.72 428.64 ;
      RECT 119.08 431.28 120.72 431.48 ;
      RECT 120.56 430.36 120.72 431.48 ;
      RECT 117.5 431.15 119.24 431.31 ;
      RECT 117.5 430.51 117.66 431.31 ;
      RECT 120.56 430.73 122.96 430.91 ;
      RECT 116.78 430.51 117.66 430.67 ;
      RECT 119.72 430.36 120.72 430.52 ;
      RECT 119.72 436.2 120.72 436.36 ;
      RECT 120.56 435.24 120.72 436.36 ;
      RECT 116.78 436.05 117.66 436.21 ;
      RECT 117.5 435.41 117.66 436.21 ;
      RECT 120.56 435.81 122.96 435.99 ;
      RECT 117.5 435.41 119.24 435.57 ;
      RECT 119.08 435.24 120.72 435.44 ;
      RECT 119.08 438.08 120.72 438.28 ;
      RECT 120.56 437.16 120.72 438.28 ;
      RECT 117.5 437.95 119.24 438.11 ;
      RECT 117.5 437.31 117.66 438.11 ;
      RECT 120.56 437.53 122.96 437.71 ;
      RECT 116.78 437.31 117.66 437.47 ;
      RECT 119.72 437.16 120.72 437.32 ;
      RECT 119.72 443 120.72 443.16 ;
      RECT 120.56 442.04 120.72 443.16 ;
      RECT 116.78 442.85 117.66 443.01 ;
      RECT 117.5 442.21 117.66 443.01 ;
      RECT 120.56 442.61 122.96 442.79 ;
      RECT 117.5 442.21 119.24 442.37 ;
      RECT 119.08 442.04 120.72 442.24 ;
      RECT 119.08 444.88 120.72 445.08 ;
      RECT 120.56 443.96 120.72 445.08 ;
      RECT 117.5 444.75 119.24 444.91 ;
      RECT 117.5 444.11 117.66 444.91 ;
      RECT 120.56 444.33 122.96 444.51 ;
      RECT 116.78 444.11 117.66 444.27 ;
      RECT 119.72 443.96 120.72 444.12 ;
      RECT 119.72 449.8 120.72 449.96 ;
      RECT 120.56 448.84 120.72 449.96 ;
      RECT 116.78 449.65 117.66 449.81 ;
      RECT 117.5 449.01 117.66 449.81 ;
      RECT 120.56 449.41 122.96 449.59 ;
      RECT 117.5 449.01 119.24 449.17 ;
      RECT 119.08 448.84 120.72 449.04 ;
      RECT 119.08 451.68 120.72 451.88 ;
      RECT 120.56 450.76 120.72 451.88 ;
      RECT 117.5 451.55 119.24 451.71 ;
      RECT 117.5 450.91 117.66 451.71 ;
      RECT 120.56 451.13 122.96 451.31 ;
      RECT 116.78 450.91 117.66 451.07 ;
      RECT 119.72 450.76 120.72 450.92 ;
      RECT 119.72 456.6 120.72 456.76 ;
      RECT 120.56 455.64 120.72 456.76 ;
      RECT 116.78 456.45 117.66 456.61 ;
      RECT 117.5 455.81 117.66 456.61 ;
      RECT 120.56 456.21 122.96 456.39 ;
      RECT 117.5 455.81 119.24 455.97 ;
      RECT 119.08 455.64 120.72 455.84 ;
      RECT 119.08 458.48 120.72 458.68 ;
      RECT 120.56 457.56 120.72 458.68 ;
      RECT 117.5 458.35 119.24 458.51 ;
      RECT 117.5 457.71 117.66 458.51 ;
      RECT 120.56 457.93 122.96 458.11 ;
      RECT 116.78 457.71 117.66 457.87 ;
      RECT 119.72 457.56 120.72 457.72 ;
      RECT 119.72 463.4 120.72 463.56 ;
      RECT 120.56 462.44 120.72 463.56 ;
      RECT 116.78 463.25 117.66 463.41 ;
      RECT 117.5 462.61 117.66 463.41 ;
      RECT 120.56 463.01 122.96 463.19 ;
      RECT 117.5 462.61 119.24 462.77 ;
      RECT 119.08 462.44 120.72 462.64 ;
      RECT 119.08 465.28 120.72 465.48 ;
      RECT 120.56 464.36 120.72 465.48 ;
      RECT 117.5 465.15 119.24 465.31 ;
      RECT 117.5 464.51 117.66 465.31 ;
      RECT 120.56 464.73 122.96 464.91 ;
      RECT 116.78 464.51 117.66 464.67 ;
      RECT 119.72 464.36 120.72 464.52 ;
      RECT 119.72 470.2 120.72 470.36 ;
      RECT 120.56 469.24 120.72 470.36 ;
      RECT 116.78 470.05 117.66 470.21 ;
      RECT 117.5 469.41 117.66 470.21 ;
      RECT 120.56 469.81 122.96 469.99 ;
      RECT 117.5 469.41 119.24 469.57 ;
      RECT 119.08 469.24 120.72 469.44 ;
      RECT 119.08 472.08 120.72 472.28 ;
      RECT 120.56 471.16 120.72 472.28 ;
      RECT 117.5 471.95 119.24 472.11 ;
      RECT 117.5 471.31 117.66 472.11 ;
      RECT 120.56 471.53 122.96 471.71 ;
      RECT 116.78 471.31 117.66 471.47 ;
      RECT 119.72 471.16 120.72 471.32 ;
      RECT 119.72 477 120.72 477.16 ;
      RECT 120.56 476.04 120.72 477.16 ;
      RECT 116.78 476.85 117.66 477.01 ;
      RECT 117.5 476.21 117.66 477.01 ;
      RECT 120.56 476.61 122.96 476.79 ;
      RECT 117.5 476.21 119.24 476.37 ;
      RECT 119.08 476.04 120.72 476.24 ;
      RECT 119.08 478.88 120.72 479.08 ;
      RECT 120.56 477.96 120.72 479.08 ;
      RECT 117.5 478.75 119.24 478.91 ;
      RECT 117.5 478.11 117.66 478.91 ;
      RECT 120.56 478.33 122.96 478.51 ;
      RECT 116.78 478.11 117.66 478.27 ;
      RECT 119.72 477.96 120.72 478.12 ;
      RECT 119.72 483.8 120.72 483.96 ;
      RECT 120.56 482.84 120.72 483.96 ;
      RECT 116.78 483.65 117.66 483.81 ;
      RECT 117.5 483.01 117.66 483.81 ;
      RECT 120.56 483.41 122.96 483.59 ;
      RECT 117.5 483.01 119.24 483.17 ;
      RECT 119.08 482.84 120.72 483.04 ;
      RECT 119.08 485.68 120.72 485.88 ;
      RECT 120.56 484.76 120.72 485.88 ;
      RECT 117.5 485.55 119.24 485.71 ;
      RECT 117.5 484.91 117.66 485.71 ;
      RECT 120.56 485.13 122.96 485.31 ;
      RECT 116.78 484.91 117.66 485.07 ;
      RECT 119.72 484.76 120.72 484.92 ;
      RECT 119.72 490.6 120.72 490.76 ;
      RECT 120.56 489.64 120.72 490.76 ;
      RECT 116.78 490.45 117.66 490.61 ;
      RECT 117.5 489.81 117.66 490.61 ;
      RECT 120.56 490.21 122.96 490.39 ;
      RECT 117.5 489.81 119.24 489.97 ;
      RECT 119.08 489.64 120.72 489.84 ;
      RECT 119.08 492.48 120.72 492.68 ;
      RECT 120.56 491.56 120.72 492.68 ;
      RECT 117.5 492.35 119.24 492.51 ;
      RECT 117.5 491.71 117.66 492.51 ;
      RECT 120.56 491.93 122.96 492.11 ;
      RECT 116.78 491.71 117.66 491.87 ;
      RECT 119.72 491.56 120.72 491.72 ;
      RECT 119.72 497.4 120.72 497.56 ;
      RECT 120.56 496.44 120.72 497.56 ;
      RECT 116.78 497.25 117.66 497.41 ;
      RECT 117.5 496.61 117.66 497.41 ;
      RECT 120.56 497.01 122.96 497.19 ;
      RECT 117.5 496.61 119.24 496.77 ;
      RECT 119.08 496.44 120.72 496.64 ;
      RECT 119.08 499.28 120.72 499.48 ;
      RECT 120.56 498.36 120.72 499.48 ;
      RECT 117.5 499.15 119.24 499.31 ;
      RECT 117.5 498.51 117.66 499.31 ;
      RECT 120.56 498.73 122.96 498.91 ;
      RECT 116.78 498.51 117.66 498.67 ;
      RECT 119.72 498.36 120.72 498.52 ;
      RECT 119.72 504.2 120.72 504.36 ;
      RECT 120.56 503.24 120.72 504.36 ;
      RECT 116.78 504.05 117.66 504.21 ;
      RECT 117.5 503.41 117.66 504.21 ;
      RECT 120.56 503.81 122.96 503.99 ;
      RECT 117.5 503.41 119.24 503.57 ;
      RECT 119.08 503.24 120.72 503.44 ;
      RECT 121.47 12.34 121.75 12.62 ;
      RECT 120.55 12.34 120.83 12.62 ;
      RECT 117.99 12.34 118.27 12.62 ;
      RECT 117.07 12.34 117.35 12.62 ;
      RECT 114.67 12.34 114.95 12.62 ;
      RECT 113.75 12.34 114.03 12.62 ;
      RECT 121.59 11.75 121.75 12.62 ;
      RECT 120.55 11.75 120.71 12.62 ;
      RECT 118.11 11.75 118.27 12.62 ;
      RECT 117.07 11.75 117.23 12.62 ;
      RECT 114.79 11.75 114.95 12.62 ;
      RECT 113.75 11.75 113.91 12.62 ;
      RECT 122.73 8.38 122.89 12.03 ;
      RECT 121.63 9.02 121.79 12.03 ;
      RECT 120.43 9.02 120.59 12.03 ;
      RECT 119.33 8.38 119.49 12.03 ;
      RECT 118.23 9.02 118.39 12.03 ;
      RECT 117.03 9.02 117.19 12.03 ;
      RECT 115.93 8.38 116.09 12.03 ;
      RECT 114.83 9.02 114.99 12.03 ;
      RECT 113.63 9.02 113.79 12.03 ;
      RECT 112.53 8.38 112.69 12.03 ;
      RECT 112.53 9.02 122.89 9.3 ;
      RECT 122.05 8.38 122.29 9.3 ;
      RECT 121.37 8.38 121.61 9.3 ;
      RECT 120.62 8.38 120.86 9.3 ;
      RECT 119.93 8.38 120.17 9.3 ;
      RECT 118.65 8.38 118.89 9.3 ;
      RECT 117.96 8.38 118.2 9.3 ;
      RECT 117.21 8.38 117.45 9.3 ;
      RECT 116.53 8.38 116.77 9.3 ;
      RECT 115.25 8.38 115.49 9.3 ;
      RECT 114.57 8.38 114.81 9.3 ;
      RECT 113.82 8.38 114.06 9.3 ;
      RECT 113.13 8.38 113.37 9.3 ;
      RECT 119.4 70.41 120.4 70.6 ;
      RECT 119.4 69.48 119.56 70.6 ;
      RECT 118.49 69.48 122.66 69.64 ;
      RECT 119.4 77.21 120.4 77.4 ;
      RECT 119.4 75.32 119.56 77.4 ;
      RECT 118.49 76.28 122.66 76.44 ;
      RECT 119.4 75.32 120.4 75.51 ;
      RECT 119.4 84.01 120.4 84.2 ;
      RECT 119.4 82.12 119.56 84.2 ;
      RECT 118.49 83.08 122.66 83.24 ;
      RECT 119.4 82.12 120.4 82.31 ;
      RECT 119.4 90.81 120.4 91 ;
      RECT 119.4 88.92 119.56 91 ;
      RECT 118.49 89.88 122.66 90.04 ;
      RECT 119.4 88.92 120.4 89.11 ;
      RECT 119.4 97.61 120.4 97.8 ;
      RECT 119.4 95.72 119.56 97.8 ;
      RECT 118.49 96.68 122.66 96.84 ;
      RECT 119.4 95.72 120.4 95.91 ;
      RECT 119.4 104.41 120.4 104.6 ;
      RECT 119.4 102.52 119.56 104.6 ;
      RECT 118.49 103.48 122.66 103.64 ;
      RECT 119.4 102.52 120.4 102.71 ;
      RECT 119.4 111.21 120.4 111.4 ;
      RECT 119.4 109.32 119.56 111.4 ;
      RECT 118.49 110.28 122.66 110.44 ;
      RECT 119.4 109.32 120.4 109.51 ;
      RECT 119.4 118.01 120.4 118.2 ;
      RECT 119.4 116.12 119.56 118.2 ;
      RECT 118.49 117.08 122.66 117.24 ;
      RECT 119.4 116.12 120.4 116.31 ;
      RECT 119.4 124.81 120.4 125 ;
      RECT 119.4 122.92 119.56 125 ;
      RECT 118.49 123.88 122.66 124.04 ;
      RECT 119.4 122.92 120.4 123.11 ;
      RECT 119.4 131.61 120.4 131.8 ;
      RECT 119.4 129.72 119.56 131.8 ;
      RECT 118.49 130.68 122.66 130.84 ;
      RECT 119.4 129.72 120.4 129.91 ;
      RECT 119.4 138.41 120.4 138.6 ;
      RECT 119.4 136.52 119.56 138.6 ;
      RECT 118.49 137.48 122.66 137.64 ;
      RECT 119.4 136.52 120.4 136.71 ;
      RECT 119.4 145.21 120.4 145.4 ;
      RECT 119.4 143.32 119.56 145.4 ;
      RECT 118.49 144.28 122.66 144.44 ;
      RECT 119.4 143.32 120.4 143.51 ;
      RECT 119.4 152.01 120.4 152.2 ;
      RECT 119.4 150.12 119.56 152.2 ;
      RECT 118.49 151.08 122.66 151.24 ;
      RECT 119.4 150.12 120.4 150.31 ;
      RECT 119.4 158.81 120.4 159 ;
      RECT 119.4 156.92 119.56 159 ;
      RECT 118.49 157.88 122.66 158.04 ;
      RECT 119.4 156.92 120.4 157.11 ;
      RECT 119.4 165.61 120.4 165.8 ;
      RECT 119.4 163.72 119.56 165.8 ;
      RECT 118.49 164.68 122.66 164.84 ;
      RECT 119.4 163.72 120.4 163.91 ;
      RECT 119.4 172.41 120.4 172.6 ;
      RECT 119.4 170.52 119.56 172.6 ;
      RECT 118.49 171.48 122.66 171.64 ;
      RECT 119.4 170.52 120.4 170.71 ;
      RECT 119.4 179.21 120.4 179.4 ;
      RECT 119.4 177.32 119.56 179.4 ;
      RECT 118.49 178.28 122.66 178.44 ;
      RECT 119.4 177.32 120.4 177.51 ;
      RECT 119.4 186.01 120.4 186.2 ;
      RECT 119.4 184.12 119.56 186.2 ;
      RECT 118.49 185.08 122.66 185.24 ;
      RECT 119.4 184.12 120.4 184.31 ;
      RECT 119.4 192.81 120.4 193 ;
      RECT 119.4 190.92 119.56 193 ;
      RECT 118.49 191.88 122.66 192.04 ;
      RECT 119.4 190.92 120.4 191.11 ;
      RECT 119.4 199.61 120.4 199.8 ;
      RECT 119.4 197.72 119.56 199.8 ;
      RECT 118.49 198.68 122.66 198.84 ;
      RECT 119.4 197.72 120.4 197.91 ;
      RECT 119.4 206.41 120.4 206.6 ;
      RECT 119.4 204.52 119.56 206.6 ;
      RECT 118.49 205.48 122.66 205.64 ;
      RECT 119.4 204.52 120.4 204.71 ;
      RECT 119.4 213.21 120.4 213.4 ;
      RECT 119.4 211.32 119.56 213.4 ;
      RECT 118.49 212.28 122.66 212.44 ;
      RECT 119.4 211.32 120.4 211.51 ;
      RECT 119.4 220.01 120.4 220.2 ;
      RECT 119.4 218.12 119.56 220.2 ;
      RECT 118.49 219.08 122.66 219.24 ;
      RECT 119.4 218.12 120.4 218.31 ;
      RECT 119.4 226.81 120.4 227 ;
      RECT 119.4 224.92 119.56 227 ;
      RECT 118.49 225.88 122.66 226.04 ;
      RECT 119.4 224.92 120.4 225.11 ;
      RECT 119.4 233.61 120.4 233.8 ;
      RECT 119.4 231.72 119.56 233.8 ;
      RECT 118.49 232.68 122.66 232.84 ;
      RECT 119.4 231.72 120.4 231.91 ;
      RECT 119.4 240.41 120.4 240.6 ;
      RECT 119.4 238.52 119.56 240.6 ;
      RECT 118.49 239.48 122.66 239.64 ;
      RECT 119.4 238.52 120.4 238.71 ;
      RECT 119.4 247.21 120.4 247.4 ;
      RECT 119.4 245.32 119.56 247.4 ;
      RECT 118.49 246.28 122.66 246.44 ;
      RECT 119.4 245.32 120.4 245.51 ;
      RECT 119.4 254.01 120.4 254.2 ;
      RECT 119.4 252.12 119.56 254.2 ;
      RECT 118.49 253.08 122.66 253.24 ;
      RECT 119.4 252.12 120.4 252.31 ;
      RECT 119.4 260.81 120.4 261 ;
      RECT 119.4 258.92 119.56 261 ;
      RECT 118.49 259.88 122.66 260.04 ;
      RECT 119.4 258.92 120.4 259.11 ;
      RECT 119.4 267.61 120.4 267.8 ;
      RECT 119.4 265.72 119.56 267.8 ;
      RECT 118.49 266.68 122.66 266.84 ;
      RECT 119.4 265.72 120.4 265.91 ;
      RECT 119.4 274.41 120.4 274.6 ;
      RECT 119.4 272.52 119.56 274.6 ;
      RECT 118.49 273.48 122.66 273.64 ;
      RECT 119.4 272.52 120.4 272.71 ;
      RECT 119.4 281.21 120.4 281.4 ;
      RECT 119.4 279.32 119.56 281.4 ;
      RECT 118.49 280.28 122.66 280.44 ;
      RECT 119.4 279.32 120.4 279.51 ;
      RECT 119.4 288.01 120.4 288.2 ;
      RECT 119.4 286.12 119.56 288.2 ;
      RECT 118.49 287.08 122.66 287.24 ;
      RECT 119.4 286.12 120.4 286.31 ;
      RECT 119.4 294.81 120.4 295 ;
      RECT 119.4 292.92 119.56 295 ;
      RECT 118.49 293.88 122.66 294.04 ;
      RECT 119.4 292.92 120.4 293.11 ;
      RECT 119.4 301.61 120.4 301.8 ;
      RECT 119.4 299.72 119.56 301.8 ;
      RECT 118.49 300.68 122.66 300.84 ;
      RECT 119.4 299.72 120.4 299.91 ;
      RECT 119.4 308.41 120.4 308.6 ;
      RECT 119.4 306.52 119.56 308.6 ;
      RECT 118.49 307.48 122.66 307.64 ;
      RECT 119.4 306.52 120.4 306.71 ;
      RECT 119.4 315.21 120.4 315.4 ;
      RECT 119.4 313.32 119.56 315.4 ;
      RECT 118.49 314.28 122.66 314.44 ;
      RECT 119.4 313.32 120.4 313.51 ;
      RECT 119.4 322.01 120.4 322.2 ;
      RECT 119.4 320.12 119.56 322.2 ;
      RECT 118.49 321.08 122.66 321.24 ;
      RECT 119.4 320.12 120.4 320.31 ;
      RECT 119.4 328.81 120.4 329 ;
      RECT 119.4 326.92 119.56 329 ;
      RECT 118.49 327.88 122.66 328.04 ;
      RECT 119.4 326.92 120.4 327.11 ;
      RECT 119.4 335.61 120.4 335.8 ;
      RECT 119.4 333.72 119.56 335.8 ;
      RECT 118.49 334.68 122.66 334.84 ;
      RECT 119.4 333.72 120.4 333.91 ;
      RECT 119.4 342.41 120.4 342.6 ;
      RECT 119.4 340.52 119.56 342.6 ;
      RECT 118.49 341.48 122.66 341.64 ;
      RECT 119.4 340.52 120.4 340.71 ;
      RECT 119.4 349.21 120.4 349.4 ;
      RECT 119.4 347.32 119.56 349.4 ;
      RECT 118.49 348.28 122.66 348.44 ;
      RECT 119.4 347.32 120.4 347.51 ;
      RECT 119.4 356.01 120.4 356.2 ;
      RECT 119.4 354.12 119.56 356.2 ;
      RECT 118.49 355.08 122.66 355.24 ;
      RECT 119.4 354.12 120.4 354.31 ;
      RECT 119.4 362.81 120.4 363 ;
      RECT 119.4 360.92 119.56 363 ;
      RECT 118.49 361.88 122.66 362.04 ;
      RECT 119.4 360.92 120.4 361.11 ;
      RECT 119.4 369.61 120.4 369.8 ;
      RECT 119.4 367.72 119.56 369.8 ;
      RECT 118.49 368.68 122.66 368.84 ;
      RECT 119.4 367.72 120.4 367.91 ;
      RECT 119.4 376.41 120.4 376.6 ;
      RECT 119.4 374.52 119.56 376.6 ;
      RECT 118.49 375.48 122.66 375.64 ;
      RECT 119.4 374.52 120.4 374.71 ;
      RECT 119.4 383.21 120.4 383.4 ;
      RECT 119.4 381.32 119.56 383.4 ;
      RECT 118.49 382.28 122.66 382.44 ;
      RECT 119.4 381.32 120.4 381.51 ;
      RECT 119.4 390.01 120.4 390.2 ;
      RECT 119.4 388.12 119.56 390.2 ;
      RECT 118.49 389.08 122.66 389.24 ;
      RECT 119.4 388.12 120.4 388.31 ;
      RECT 119.4 396.81 120.4 397 ;
      RECT 119.4 394.92 119.56 397 ;
      RECT 118.49 395.88 122.66 396.04 ;
      RECT 119.4 394.92 120.4 395.11 ;
      RECT 119.4 403.61 120.4 403.8 ;
      RECT 119.4 401.72 119.56 403.8 ;
      RECT 118.49 402.68 122.66 402.84 ;
      RECT 119.4 401.72 120.4 401.91 ;
      RECT 119.4 410.41 120.4 410.6 ;
      RECT 119.4 408.52 119.56 410.6 ;
      RECT 118.49 409.48 122.66 409.64 ;
      RECT 119.4 408.52 120.4 408.71 ;
      RECT 119.4 417.21 120.4 417.4 ;
      RECT 119.4 415.32 119.56 417.4 ;
      RECT 118.49 416.28 122.66 416.44 ;
      RECT 119.4 415.32 120.4 415.51 ;
      RECT 119.4 424.01 120.4 424.2 ;
      RECT 119.4 422.12 119.56 424.2 ;
      RECT 118.49 423.08 122.66 423.24 ;
      RECT 119.4 422.12 120.4 422.31 ;
      RECT 119.4 430.81 120.4 431 ;
      RECT 119.4 428.92 119.56 431 ;
      RECT 118.49 429.88 122.66 430.04 ;
      RECT 119.4 428.92 120.4 429.11 ;
      RECT 119.4 437.61 120.4 437.8 ;
      RECT 119.4 435.72 119.56 437.8 ;
      RECT 118.49 436.68 122.66 436.84 ;
      RECT 119.4 435.72 120.4 435.91 ;
      RECT 119.4 444.41 120.4 444.6 ;
      RECT 119.4 442.52 119.56 444.6 ;
      RECT 118.49 443.48 122.66 443.64 ;
      RECT 119.4 442.52 120.4 442.71 ;
      RECT 119.4 451.21 120.4 451.4 ;
      RECT 119.4 449.32 119.56 451.4 ;
      RECT 118.49 450.28 122.66 450.44 ;
      RECT 119.4 449.32 120.4 449.51 ;
      RECT 119.4 458.01 120.4 458.2 ;
      RECT 119.4 456.12 119.56 458.2 ;
      RECT 118.49 457.08 122.66 457.24 ;
      RECT 119.4 456.12 120.4 456.31 ;
      RECT 119.4 464.81 120.4 465 ;
      RECT 119.4 462.92 119.56 465 ;
      RECT 118.49 463.88 122.66 464.04 ;
      RECT 119.4 462.92 120.4 463.11 ;
      RECT 119.4 471.61 120.4 471.8 ;
      RECT 119.4 469.72 119.56 471.8 ;
      RECT 118.49 470.68 122.66 470.84 ;
      RECT 119.4 469.72 120.4 469.91 ;
      RECT 119.4 478.41 120.4 478.6 ;
      RECT 119.4 476.52 119.56 478.6 ;
      RECT 118.49 477.48 122.66 477.64 ;
      RECT 119.4 476.52 120.4 476.71 ;
      RECT 119.4 485.21 120.4 485.4 ;
      RECT 119.4 483.32 119.56 485.4 ;
      RECT 118.49 484.28 122.66 484.44 ;
      RECT 119.4 483.32 120.4 483.51 ;
      RECT 119.4 492.01 120.4 492.2 ;
      RECT 119.4 490.12 119.56 492.2 ;
      RECT 118.49 491.08 122.66 491.24 ;
      RECT 119.4 490.12 120.4 490.31 ;
      RECT 119.4 498.81 120.4 499 ;
      RECT 119.4 496.92 119.56 499 ;
      RECT 118.49 497.88 122.66 498.04 ;
      RECT 119.4 496.92 120.4 497.11 ;
      RECT 119.4 73.84 120.4 74 ;
      RECT 119.4 71.92 119.56 74 ;
      RECT 118.49 72.88 122.58 73.04 ;
      RECT 119.4 71.92 120.4 72.08 ;
      RECT 119.4 80.64 120.4 80.8 ;
      RECT 119.4 78.72 119.56 80.8 ;
      RECT 118.49 79.68 122.58 79.84 ;
      RECT 119.4 78.72 120.4 78.88 ;
      RECT 119.4 87.44 120.4 87.6 ;
      RECT 119.4 85.52 119.56 87.6 ;
      RECT 118.49 86.48 122.58 86.64 ;
      RECT 119.4 85.52 120.4 85.68 ;
      RECT 119.4 94.24 120.4 94.4 ;
      RECT 119.4 92.32 119.56 94.4 ;
      RECT 118.49 93.28 122.58 93.44 ;
      RECT 119.4 92.32 120.4 92.48 ;
      RECT 119.4 101.04 120.4 101.2 ;
      RECT 119.4 99.12 119.56 101.2 ;
      RECT 118.49 100.08 122.58 100.24 ;
      RECT 119.4 99.12 120.4 99.28 ;
      RECT 119.4 107.84 120.4 108 ;
      RECT 119.4 105.92 119.56 108 ;
      RECT 118.49 106.88 122.58 107.04 ;
      RECT 119.4 105.92 120.4 106.08 ;
      RECT 119.4 114.64 120.4 114.8 ;
      RECT 119.4 112.72 119.56 114.8 ;
      RECT 118.49 113.68 122.58 113.84 ;
      RECT 119.4 112.72 120.4 112.88 ;
      RECT 119.4 121.44 120.4 121.6 ;
      RECT 119.4 119.52 119.56 121.6 ;
      RECT 118.49 120.48 122.58 120.64 ;
      RECT 119.4 119.52 120.4 119.68 ;
      RECT 119.4 128.24 120.4 128.4 ;
      RECT 119.4 126.32 119.56 128.4 ;
      RECT 118.49 127.28 122.58 127.44 ;
      RECT 119.4 126.32 120.4 126.48 ;
      RECT 119.4 135.04 120.4 135.2 ;
      RECT 119.4 133.12 119.56 135.2 ;
      RECT 118.49 134.08 122.58 134.24 ;
      RECT 119.4 133.12 120.4 133.28 ;
      RECT 119.4 141.84 120.4 142 ;
      RECT 119.4 139.92 119.56 142 ;
      RECT 118.49 140.88 122.58 141.04 ;
      RECT 119.4 139.92 120.4 140.08 ;
      RECT 119.4 148.64 120.4 148.8 ;
      RECT 119.4 146.72 119.56 148.8 ;
      RECT 118.49 147.68 122.58 147.84 ;
      RECT 119.4 146.72 120.4 146.88 ;
      RECT 119.4 155.44 120.4 155.6 ;
      RECT 119.4 153.52 119.56 155.6 ;
      RECT 118.49 154.48 122.58 154.64 ;
      RECT 119.4 153.52 120.4 153.68 ;
      RECT 119.4 162.24 120.4 162.4 ;
      RECT 119.4 160.32 119.56 162.4 ;
      RECT 118.49 161.28 122.58 161.44 ;
      RECT 119.4 160.32 120.4 160.48 ;
      RECT 119.4 169.04 120.4 169.2 ;
      RECT 119.4 167.12 119.56 169.2 ;
      RECT 118.49 168.08 122.58 168.24 ;
      RECT 119.4 167.12 120.4 167.28 ;
      RECT 119.4 175.84 120.4 176 ;
      RECT 119.4 173.92 119.56 176 ;
      RECT 118.49 174.88 122.58 175.04 ;
      RECT 119.4 173.92 120.4 174.08 ;
      RECT 119.4 182.64 120.4 182.8 ;
      RECT 119.4 180.72 119.56 182.8 ;
      RECT 118.49 181.68 122.58 181.84 ;
      RECT 119.4 180.72 120.4 180.88 ;
      RECT 119.4 189.44 120.4 189.6 ;
      RECT 119.4 187.52 119.56 189.6 ;
      RECT 118.49 188.48 122.58 188.64 ;
      RECT 119.4 187.52 120.4 187.68 ;
      RECT 119.4 196.24 120.4 196.4 ;
      RECT 119.4 194.32 119.56 196.4 ;
      RECT 118.49 195.28 122.58 195.44 ;
      RECT 119.4 194.32 120.4 194.48 ;
      RECT 119.4 203.04 120.4 203.2 ;
      RECT 119.4 201.12 119.56 203.2 ;
      RECT 118.49 202.08 122.58 202.24 ;
      RECT 119.4 201.12 120.4 201.28 ;
      RECT 119.4 209.84 120.4 210 ;
      RECT 119.4 207.92 119.56 210 ;
      RECT 118.49 208.88 122.58 209.04 ;
      RECT 119.4 207.92 120.4 208.08 ;
      RECT 119.4 216.64 120.4 216.8 ;
      RECT 119.4 214.72 119.56 216.8 ;
      RECT 118.49 215.68 122.58 215.84 ;
      RECT 119.4 214.72 120.4 214.88 ;
      RECT 119.4 223.44 120.4 223.6 ;
      RECT 119.4 221.52 119.56 223.6 ;
      RECT 118.49 222.48 122.58 222.64 ;
      RECT 119.4 221.52 120.4 221.68 ;
      RECT 119.4 230.24 120.4 230.4 ;
      RECT 119.4 228.32 119.56 230.4 ;
      RECT 118.49 229.28 122.58 229.44 ;
      RECT 119.4 228.32 120.4 228.48 ;
      RECT 119.4 237.04 120.4 237.2 ;
      RECT 119.4 235.12 119.56 237.2 ;
      RECT 118.49 236.08 122.58 236.24 ;
      RECT 119.4 235.12 120.4 235.28 ;
      RECT 119.4 243.84 120.4 244 ;
      RECT 119.4 241.92 119.56 244 ;
      RECT 118.49 242.88 122.58 243.04 ;
      RECT 119.4 241.92 120.4 242.08 ;
      RECT 119.4 250.64 120.4 250.8 ;
      RECT 119.4 248.72 119.56 250.8 ;
      RECT 118.49 249.68 122.58 249.84 ;
      RECT 119.4 248.72 120.4 248.88 ;
      RECT 119.4 257.44 120.4 257.6 ;
      RECT 119.4 255.52 119.56 257.6 ;
      RECT 118.49 256.48 122.58 256.64 ;
      RECT 119.4 255.52 120.4 255.68 ;
      RECT 119.4 264.24 120.4 264.4 ;
      RECT 119.4 262.32 119.56 264.4 ;
      RECT 118.49 263.28 122.58 263.44 ;
      RECT 119.4 262.32 120.4 262.48 ;
      RECT 119.4 271.04 120.4 271.2 ;
      RECT 119.4 269.12 119.56 271.2 ;
      RECT 118.49 270.08 122.58 270.24 ;
      RECT 119.4 269.12 120.4 269.28 ;
      RECT 119.4 277.84 120.4 278 ;
      RECT 119.4 275.92 119.56 278 ;
      RECT 118.49 276.88 122.58 277.04 ;
      RECT 119.4 275.92 120.4 276.08 ;
      RECT 119.4 284.64 120.4 284.8 ;
      RECT 119.4 282.72 119.56 284.8 ;
      RECT 118.49 283.68 122.58 283.84 ;
      RECT 119.4 282.72 120.4 282.88 ;
      RECT 119.4 291.44 120.4 291.6 ;
      RECT 119.4 289.52 119.56 291.6 ;
      RECT 118.49 290.48 122.58 290.64 ;
      RECT 119.4 289.52 120.4 289.68 ;
      RECT 119.4 298.24 120.4 298.4 ;
      RECT 119.4 296.32 119.56 298.4 ;
      RECT 118.49 297.28 122.58 297.44 ;
      RECT 119.4 296.32 120.4 296.48 ;
      RECT 119.4 305.04 120.4 305.2 ;
      RECT 119.4 303.12 119.56 305.2 ;
      RECT 118.49 304.08 122.58 304.24 ;
      RECT 119.4 303.12 120.4 303.28 ;
      RECT 119.4 311.84 120.4 312 ;
      RECT 119.4 309.92 119.56 312 ;
      RECT 118.49 310.88 122.58 311.04 ;
      RECT 119.4 309.92 120.4 310.08 ;
      RECT 119.4 318.64 120.4 318.8 ;
      RECT 119.4 316.72 119.56 318.8 ;
      RECT 118.49 317.68 122.58 317.84 ;
      RECT 119.4 316.72 120.4 316.88 ;
      RECT 119.4 325.44 120.4 325.6 ;
      RECT 119.4 323.52 119.56 325.6 ;
      RECT 118.49 324.48 122.58 324.64 ;
      RECT 119.4 323.52 120.4 323.68 ;
      RECT 119.4 332.24 120.4 332.4 ;
      RECT 119.4 330.32 119.56 332.4 ;
      RECT 118.49 331.28 122.58 331.44 ;
      RECT 119.4 330.32 120.4 330.48 ;
      RECT 119.4 339.04 120.4 339.2 ;
      RECT 119.4 337.12 119.56 339.2 ;
      RECT 118.49 338.08 122.58 338.24 ;
      RECT 119.4 337.12 120.4 337.28 ;
      RECT 119.4 345.84 120.4 346 ;
      RECT 119.4 343.92 119.56 346 ;
      RECT 118.49 344.88 122.58 345.04 ;
      RECT 119.4 343.92 120.4 344.08 ;
      RECT 119.4 352.64 120.4 352.8 ;
      RECT 119.4 350.72 119.56 352.8 ;
      RECT 118.49 351.68 122.58 351.84 ;
      RECT 119.4 350.72 120.4 350.88 ;
      RECT 119.4 359.44 120.4 359.6 ;
      RECT 119.4 357.52 119.56 359.6 ;
      RECT 118.49 358.48 122.58 358.64 ;
      RECT 119.4 357.52 120.4 357.68 ;
      RECT 119.4 366.24 120.4 366.4 ;
      RECT 119.4 364.32 119.56 366.4 ;
      RECT 118.49 365.28 122.58 365.44 ;
      RECT 119.4 364.32 120.4 364.48 ;
      RECT 119.4 373.04 120.4 373.2 ;
      RECT 119.4 371.12 119.56 373.2 ;
      RECT 118.49 372.08 122.58 372.24 ;
      RECT 119.4 371.12 120.4 371.28 ;
      RECT 119.4 379.84 120.4 380 ;
      RECT 119.4 377.92 119.56 380 ;
      RECT 118.49 378.88 122.58 379.04 ;
      RECT 119.4 377.92 120.4 378.08 ;
      RECT 119.4 386.64 120.4 386.8 ;
      RECT 119.4 384.72 119.56 386.8 ;
      RECT 118.49 385.68 122.58 385.84 ;
      RECT 119.4 384.72 120.4 384.88 ;
      RECT 119.4 393.44 120.4 393.6 ;
      RECT 119.4 391.52 119.56 393.6 ;
      RECT 118.49 392.48 122.58 392.64 ;
      RECT 119.4 391.52 120.4 391.68 ;
      RECT 119.4 400.24 120.4 400.4 ;
      RECT 119.4 398.32 119.56 400.4 ;
      RECT 118.49 399.28 122.58 399.44 ;
      RECT 119.4 398.32 120.4 398.48 ;
      RECT 119.4 407.04 120.4 407.2 ;
      RECT 119.4 405.12 119.56 407.2 ;
      RECT 118.49 406.08 122.58 406.24 ;
      RECT 119.4 405.12 120.4 405.28 ;
      RECT 119.4 413.84 120.4 414 ;
      RECT 119.4 411.92 119.56 414 ;
      RECT 118.49 412.88 122.58 413.04 ;
      RECT 119.4 411.92 120.4 412.08 ;
      RECT 119.4 420.64 120.4 420.8 ;
      RECT 119.4 418.72 119.56 420.8 ;
      RECT 118.49 419.68 122.58 419.84 ;
      RECT 119.4 418.72 120.4 418.88 ;
      RECT 119.4 427.44 120.4 427.6 ;
      RECT 119.4 425.52 119.56 427.6 ;
      RECT 118.49 426.48 122.58 426.64 ;
      RECT 119.4 425.52 120.4 425.68 ;
      RECT 119.4 434.24 120.4 434.4 ;
      RECT 119.4 432.32 119.56 434.4 ;
      RECT 118.49 433.28 122.58 433.44 ;
      RECT 119.4 432.32 120.4 432.48 ;
      RECT 119.4 441.04 120.4 441.2 ;
      RECT 119.4 439.12 119.56 441.2 ;
      RECT 118.49 440.08 122.58 440.24 ;
      RECT 119.4 439.12 120.4 439.28 ;
      RECT 119.4 447.84 120.4 448 ;
      RECT 119.4 445.92 119.56 448 ;
      RECT 118.49 446.88 122.58 447.04 ;
      RECT 119.4 445.92 120.4 446.08 ;
      RECT 119.4 454.64 120.4 454.8 ;
      RECT 119.4 452.72 119.56 454.8 ;
      RECT 118.49 453.68 122.58 453.84 ;
      RECT 119.4 452.72 120.4 452.88 ;
      RECT 119.4 461.44 120.4 461.6 ;
      RECT 119.4 459.52 119.56 461.6 ;
      RECT 118.49 460.48 122.58 460.64 ;
      RECT 119.4 459.52 120.4 459.68 ;
      RECT 119.4 468.24 120.4 468.4 ;
      RECT 119.4 466.32 119.56 468.4 ;
      RECT 118.49 467.28 122.58 467.44 ;
      RECT 119.4 466.32 120.4 466.48 ;
      RECT 119.4 475.04 120.4 475.2 ;
      RECT 119.4 473.12 119.56 475.2 ;
      RECT 118.49 474.08 122.58 474.24 ;
      RECT 119.4 473.12 120.4 473.28 ;
      RECT 119.4 481.84 120.4 482 ;
      RECT 119.4 479.92 119.56 482 ;
      RECT 118.49 480.88 122.58 481.04 ;
      RECT 119.4 479.92 120.4 480.08 ;
      RECT 119.4 488.64 120.4 488.8 ;
      RECT 119.4 486.72 119.56 488.8 ;
      RECT 118.49 487.68 122.58 487.84 ;
      RECT 119.4 486.72 120.4 486.88 ;
      RECT 119.4 495.44 120.4 495.6 ;
      RECT 119.4 493.52 119.56 495.6 ;
      RECT 118.49 494.48 122.58 494.64 ;
      RECT 119.4 493.52 120.4 493.68 ;
      RECT 119.4 502.24 120.4 502.4 ;
      RECT 119.4 500.32 119.56 502.4 ;
      RECT 118.49 501.28 122.58 501.44 ;
      RECT 119.4 500.32 120.4 500.48 ;
      RECT 121.95 49.6 122.11 51.7 ;
      RECT 121.95 49.6 122.55 49.76 ;
      RECT 122.39 32.06 122.55 49.76 ;
      RECT 121.73 45.9 122.55 46.06 ;
      RECT 121.73 36.23 122.55 36.39 ;
      RECT 121.95 32.06 122.55 32.22 ;
      RECT 121.95 30.54 122.11 32.22 ;
      RECT 120.45 21.06 120.61 26.28 ;
      RECT 121.41 24.37 121.57 25.98 ;
      RECT 120.45 24.37 121.77 24.53 ;
      RECT 121.61 23.67 121.77 24.53 ;
      RECT 121.41 23.67 121.77 23.83 ;
      RECT 121.41 21.7 121.57 23.83 ;
      RECT 120.39 21.06 122.27 21.22 ;
      RECT 120.39 60.83 122.27 60.99 ;
      RECT 120.45 55.81 120.61 60.99 ;
      RECT 121.41 58.22 121.57 60.35 ;
      RECT 121.41 58.22 121.77 58.38 ;
      RECT 121.61 57.25 121.77 58.38 ;
      RECT 120.45 57.25 121.77 57.41 ;
      RECT 121.41 56.13 121.57 57.41 ;
      RECT 120.05 25.79 120.29 26.07 ;
      RECT 120.13 21.94 120.29 26.07 ;
      RECT 120.01 21.94 120.29 22.18 ;
      RECT 120.07 15.28 120.23 22.18 ;
      RECT 121.99 15.28 122.15 20.88 ;
      RECT 121.03 15.28 121.19 20.88 ;
      RECT 120.07 17.14 122.15 17.3 ;
      RECT 120.07 35.91 122.15 36.07 ;
      RECT 121.99 32.85 122.15 36.07 ;
      RECT 121.03 27.43 121.19 36.07 ;
      RECT 120.07 32.85 120.23 36.07 ;
      RECT 121.03 27.43 122.09 27.59 ;
      RECT 121.93 23.41 122.09 27.59 ;
      RECT 120.93 26.14 122.09 26.3 ;
      RECT 121.89 25 122.09 26.3 ;
      RECT 120.93 25.01 121.09 26.3 ;
      RECT 120.93 21.38 121.09 23.81 ;
      RECT 121.89 21.38 122.05 23.55 ;
      RECT 120.93 21.38 122.05 21.54 ;
      RECT 120.93 60.51 122.05 60.67 ;
      RECT 121.89 58.5 122.05 60.67 ;
      RECT 121.93 55.81 122.05 60.67 ;
      RECT 120.93 58.24 121.09 60.67 ;
      RECT 121.95 54.64 122.09 58.64 ;
      RECT 121.89 55.81 122.11 57.09 ;
      RECT 121.95 54.64 122.11 57.09 ;
      RECT 120.93 55.81 121.09 57.09 ;
      RECT 120.93 55.81 122.11 55.97 ;
      RECT 121.03 54.64 122.11 54.8 ;
      RECT 121.03 46.22 121.19 54.8 ;
      RECT 121.99 46.22 122.15 49.44 ;
      RECT 120.07 46.22 120.23 49.44 ;
      RECT 120.07 46.22 122.15 46.38 ;
      RECT 121.99 61.17 122.15 66.77 ;
      RECT 121.03 61.17 121.19 66.77 ;
      RECT 120.07 59.87 120.23 66.77 ;
      RECT 120.07 64.75 122.15 64.91 ;
      RECT 120.01 59.87 120.29 60.11 ;
      RECT 120.13 56.02 120.29 60.11 ;
      RECT 120.05 56.02 120.29 56.3 ;
      RECT 121.03 10.09 121.19 14.2 ;
      RECT 121.03 12.9 122.09 13.06 ;
      RECT 121.93 12.19 122.09 13.06 ;
      RECT 121.91 41.08 122.07 45.17 ;
      RECT 121.75 41.08 122.07 41.24 ;
      RECT 121.51 14.52 121.67 16.86 ;
      RECT 121.64 13.22 121.8 14.84 ;
      RECT 121.51 31.09 121.67 35.75 ;
      RECT 121.51 32.25 121.77 32.53 ;
      RECT 119.73 26.46 121.75 26.62 ;
      RECT 119.73 25.35 119.89 26.62 ;
      RECT 119.81 22.91 119.97 25.51 ;
      RECT 119.81 56.46 119.97 59.14 ;
      RECT 119.73 55.49 119.89 56.62 ;
      RECT 119.73 55.49 121.75 55.65 ;
      RECT 121.51 49.75 121.71 51.3 ;
      RECT 121.51 46.54 121.67 51.3 ;
      RECT 120.39 55.09 121.65 55.25 ;
      RECT 120.39 49.77 120.55 55.25 ;
      RECT 119.67 49.77 120.55 49.93 ;
      RECT 119.67 32.48 119.83 49.93 ;
      RECT 119.67 45.9 120.49 46.06 ;
      RECT 119.67 36.23 120.49 36.39 ;
      RECT 119.67 32.48 120.55 32.64 ;
      RECT 120.39 27.04 120.55 32.64 ;
      RECT 120.39 27.04 121.65 27.2 ;
      RECT 120.77 45.9 121.57 46.06 ;
      RECT 121.41 44.89 121.57 46.06 ;
      RECT 121.43 38.57 121.59 45.17 ;
      RECT 120.63 38.57 120.79 45.17 ;
      RECT 120.63 38.57 121.09 38.73 ;
      RECT 120.93 36.23 121.09 38.73 ;
      RECT 120.77 36.23 121.45 36.39 ;
      RECT 120.55 32.85 120.71 35.75 ;
      RECT 120.71 31.09 120.87 33.01 ;
      RECT 120.71 49.44 120.87 51.3 ;
      RECT 120.55 46.54 120.71 49.6 ;
      RECT 120.13 12.8 120.79 13.06 ;
      RECT 120.13 12.19 120.37 13.06 ;
      RECT 120.55 14.52 120.71 16.86 ;
      RECT 120.42 13.22 120.58 14.84 ;
      RECT 120.15 41.08 120.31 45.17 ;
      RECT 120.15 41.08 120.47 41.24 ;
      RECT 119.33 17.6 119.49 23.81 ;
      RECT 118.85 22.38 119.97 22.54 ;
      RECT 119.33 58.24 119.49 64 ;
      RECT 118.85 59.51 119.97 59.67 ;
      RECT 119.75 27.37 119.91 31.49 ;
      RECT 118.91 27.37 119.07 31.49 ;
      RECT 118.91 27.37 119.91 27.53 ;
      RECT 119.33 24.64 119.49 27.53 ;
      RECT 119.33 54.16 119.49 57.42 ;
      RECT 118.91 54.16 119.91 54.88 ;
      RECT 119.75 50.8 119.91 54.88 ;
      RECT 118.91 50.8 119.07 54.88 ;
      RECT 118.23 70.31 118.95 70.56 ;
      RECT 118.79 69.8 118.95 70.56 ;
      RECT 117.82 70.31 118.95 70.47 ;
      RECT 118.79 69.8 119.24 69.96 ;
      RECT 118.79 72.56 119.24 72.72 ;
      RECT 118.79 71.95 118.95 72.72 ;
      RECT 117.82 72.15 118.95 72.31 ;
      RECT 118.23 71.95 118.95 72.31 ;
      RECT 118.23 73.61 118.95 73.97 ;
      RECT 118.79 73.2 118.95 73.97 ;
      RECT 117.82 73.61 118.95 73.77 ;
      RECT 118.79 73.2 119.24 73.36 ;
      RECT 118.79 75.96 119.24 76.12 ;
      RECT 118.79 75.36 118.95 76.12 ;
      RECT 117.82 75.45 118.95 75.61 ;
      RECT 118.23 75.36 118.95 75.61 ;
      RECT 118.23 77.11 118.95 77.36 ;
      RECT 118.79 76.6 118.95 77.36 ;
      RECT 117.82 77.11 118.95 77.27 ;
      RECT 118.79 76.6 119.24 76.76 ;
      RECT 118.79 79.36 119.24 79.52 ;
      RECT 118.79 78.75 118.95 79.52 ;
      RECT 117.82 78.95 118.95 79.11 ;
      RECT 118.23 78.75 118.95 79.11 ;
      RECT 118.23 80.41 118.95 80.77 ;
      RECT 118.79 80 118.95 80.77 ;
      RECT 117.82 80.41 118.95 80.57 ;
      RECT 118.79 80 119.24 80.16 ;
      RECT 118.79 82.76 119.24 82.92 ;
      RECT 118.79 82.16 118.95 82.92 ;
      RECT 117.82 82.25 118.95 82.41 ;
      RECT 118.23 82.16 118.95 82.41 ;
      RECT 118.23 83.91 118.95 84.16 ;
      RECT 118.79 83.4 118.95 84.16 ;
      RECT 117.82 83.91 118.95 84.07 ;
      RECT 118.79 83.4 119.24 83.56 ;
      RECT 118.79 86.16 119.24 86.32 ;
      RECT 118.79 85.55 118.95 86.32 ;
      RECT 117.82 85.75 118.95 85.91 ;
      RECT 118.23 85.55 118.95 85.91 ;
      RECT 118.23 87.21 118.95 87.57 ;
      RECT 118.79 86.8 118.95 87.57 ;
      RECT 117.82 87.21 118.95 87.37 ;
      RECT 118.79 86.8 119.24 86.96 ;
      RECT 118.79 89.56 119.24 89.72 ;
      RECT 118.79 88.96 118.95 89.72 ;
      RECT 117.82 89.05 118.95 89.21 ;
      RECT 118.23 88.96 118.95 89.21 ;
      RECT 118.23 90.71 118.95 90.96 ;
      RECT 118.79 90.2 118.95 90.96 ;
      RECT 117.82 90.71 118.95 90.87 ;
      RECT 118.79 90.2 119.24 90.36 ;
      RECT 118.79 92.96 119.24 93.12 ;
      RECT 118.79 92.35 118.95 93.12 ;
      RECT 117.82 92.55 118.95 92.71 ;
      RECT 118.23 92.35 118.95 92.71 ;
      RECT 118.23 94.01 118.95 94.37 ;
      RECT 118.79 93.6 118.95 94.37 ;
      RECT 117.82 94.01 118.95 94.17 ;
      RECT 118.79 93.6 119.24 93.76 ;
      RECT 118.79 96.36 119.24 96.52 ;
      RECT 118.79 95.76 118.95 96.52 ;
      RECT 117.82 95.85 118.95 96.01 ;
      RECT 118.23 95.76 118.95 96.01 ;
      RECT 118.23 97.51 118.95 97.76 ;
      RECT 118.79 97 118.95 97.76 ;
      RECT 117.82 97.51 118.95 97.67 ;
      RECT 118.79 97 119.24 97.16 ;
      RECT 118.79 99.76 119.24 99.92 ;
      RECT 118.79 99.15 118.95 99.92 ;
      RECT 117.82 99.35 118.95 99.51 ;
      RECT 118.23 99.15 118.95 99.51 ;
      RECT 118.23 100.81 118.95 101.17 ;
      RECT 118.79 100.4 118.95 101.17 ;
      RECT 117.82 100.81 118.95 100.97 ;
      RECT 118.79 100.4 119.24 100.56 ;
      RECT 118.79 103.16 119.24 103.32 ;
      RECT 118.79 102.56 118.95 103.32 ;
      RECT 117.82 102.65 118.95 102.81 ;
      RECT 118.23 102.56 118.95 102.81 ;
      RECT 118.23 104.31 118.95 104.56 ;
      RECT 118.79 103.8 118.95 104.56 ;
      RECT 117.82 104.31 118.95 104.47 ;
      RECT 118.79 103.8 119.24 103.96 ;
      RECT 118.79 106.56 119.24 106.72 ;
      RECT 118.79 105.95 118.95 106.72 ;
      RECT 117.82 106.15 118.95 106.31 ;
      RECT 118.23 105.95 118.95 106.31 ;
      RECT 118.23 107.61 118.95 107.97 ;
      RECT 118.79 107.2 118.95 107.97 ;
      RECT 117.82 107.61 118.95 107.77 ;
      RECT 118.79 107.2 119.24 107.36 ;
      RECT 118.79 109.96 119.24 110.12 ;
      RECT 118.79 109.36 118.95 110.12 ;
      RECT 117.82 109.45 118.95 109.61 ;
      RECT 118.23 109.36 118.95 109.61 ;
      RECT 118.23 111.11 118.95 111.36 ;
      RECT 118.79 110.6 118.95 111.36 ;
      RECT 117.82 111.11 118.95 111.27 ;
      RECT 118.79 110.6 119.24 110.76 ;
      RECT 118.79 113.36 119.24 113.52 ;
      RECT 118.79 112.75 118.95 113.52 ;
      RECT 117.82 112.95 118.95 113.11 ;
      RECT 118.23 112.75 118.95 113.11 ;
      RECT 118.23 114.41 118.95 114.77 ;
      RECT 118.79 114 118.95 114.77 ;
      RECT 117.82 114.41 118.95 114.57 ;
      RECT 118.79 114 119.24 114.16 ;
      RECT 118.79 116.76 119.24 116.92 ;
      RECT 118.79 116.16 118.95 116.92 ;
      RECT 117.82 116.25 118.95 116.41 ;
      RECT 118.23 116.16 118.95 116.41 ;
      RECT 118.23 117.91 118.95 118.16 ;
      RECT 118.79 117.4 118.95 118.16 ;
      RECT 117.82 117.91 118.95 118.07 ;
      RECT 118.79 117.4 119.24 117.56 ;
      RECT 118.79 120.16 119.24 120.32 ;
      RECT 118.79 119.55 118.95 120.32 ;
      RECT 117.82 119.75 118.95 119.91 ;
      RECT 118.23 119.55 118.95 119.91 ;
      RECT 118.23 121.21 118.95 121.57 ;
      RECT 118.79 120.8 118.95 121.57 ;
      RECT 117.82 121.21 118.95 121.37 ;
      RECT 118.79 120.8 119.24 120.96 ;
      RECT 118.79 123.56 119.24 123.72 ;
      RECT 118.79 122.96 118.95 123.72 ;
      RECT 117.82 123.05 118.95 123.21 ;
      RECT 118.23 122.96 118.95 123.21 ;
      RECT 118.23 124.71 118.95 124.96 ;
      RECT 118.79 124.2 118.95 124.96 ;
      RECT 117.82 124.71 118.95 124.87 ;
      RECT 118.79 124.2 119.24 124.36 ;
      RECT 118.79 126.96 119.24 127.12 ;
      RECT 118.79 126.35 118.95 127.12 ;
      RECT 117.82 126.55 118.95 126.71 ;
      RECT 118.23 126.35 118.95 126.71 ;
      RECT 118.23 128.01 118.95 128.37 ;
      RECT 118.79 127.6 118.95 128.37 ;
      RECT 117.82 128.01 118.95 128.17 ;
      RECT 118.79 127.6 119.24 127.76 ;
      RECT 118.79 130.36 119.24 130.52 ;
      RECT 118.79 129.76 118.95 130.52 ;
      RECT 117.82 129.85 118.95 130.01 ;
      RECT 118.23 129.76 118.95 130.01 ;
      RECT 118.23 131.51 118.95 131.76 ;
      RECT 118.79 131 118.95 131.76 ;
      RECT 117.82 131.51 118.95 131.67 ;
      RECT 118.79 131 119.24 131.16 ;
      RECT 118.79 133.76 119.24 133.92 ;
      RECT 118.79 133.15 118.95 133.92 ;
      RECT 117.82 133.35 118.95 133.51 ;
      RECT 118.23 133.15 118.95 133.51 ;
      RECT 118.23 134.81 118.95 135.17 ;
      RECT 118.79 134.4 118.95 135.17 ;
      RECT 117.82 134.81 118.95 134.97 ;
      RECT 118.79 134.4 119.24 134.56 ;
      RECT 118.79 137.16 119.24 137.32 ;
      RECT 118.79 136.56 118.95 137.32 ;
      RECT 117.82 136.65 118.95 136.81 ;
      RECT 118.23 136.56 118.95 136.81 ;
      RECT 118.23 138.31 118.95 138.56 ;
      RECT 118.79 137.8 118.95 138.56 ;
      RECT 117.82 138.31 118.95 138.47 ;
      RECT 118.79 137.8 119.24 137.96 ;
      RECT 118.79 140.56 119.24 140.72 ;
      RECT 118.79 139.95 118.95 140.72 ;
      RECT 117.82 140.15 118.95 140.31 ;
      RECT 118.23 139.95 118.95 140.31 ;
      RECT 118.23 141.61 118.95 141.97 ;
      RECT 118.79 141.2 118.95 141.97 ;
      RECT 117.82 141.61 118.95 141.77 ;
      RECT 118.79 141.2 119.24 141.36 ;
      RECT 118.79 143.96 119.24 144.12 ;
      RECT 118.79 143.36 118.95 144.12 ;
      RECT 117.82 143.45 118.95 143.61 ;
      RECT 118.23 143.36 118.95 143.61 ;
      RECT 118.23 145.11 118.95 145.36 ;
      RECT 118.79 144.6 118.95 145.36 ;
      RECT 117.82 145.11 118.95 145.27 ;
      RECT 118.79 144.6 119.24 144.76 ;
      RECT 118.79 147.36 119.24 147.52 ;
      RECT 118.79 146.75 118.95 147.52 ;
      RECT 117.82 146.95 118.95 147.11 ;
      RECT 118.23 146.75 118.95 147.11 ;
      RECT 118.23 148.41 118.95 148.77 ;
      RECT 118.79 148 118.95 148.77 ;
      RECT 117.82 148.41 118.95 148.57 ;
      RECT 118.79 148 119.24 148.16 ;
      RECT 118.79 150.76 119.24 150.92 ;
      RECT 118.79 150.16 118.95 150.92 ;
      RECT 117.82 150.25 118.95 150.41 ;
      RECT 118.23 150.16 118.95 150.41 ;
      RECT 118.23 151.91 118.95 152.16 ;
      RECT 118.79 151.4 118.95 152.16 ;
      RECT 117.82 151.91 118.95 152.07 ;
      RECT 118.79 151.4 119.24 151.56 ;
      RECT 118.79 154.16 119.24 154.32 ;
      RECT 118.79 153.55 118.95 154.32 ;
      RECT 117.82 153.75 118.95 153.91 ;
      RECT 118.23 153.55 118.95 153.91 ;
      RECT 118.23 155.21 118.95 155.57 ;
      RECT 118.79 154.8 118.95 155.57 ;
      RECT 117.82 155.21 118.95 155.37 ;
      RECT 118.79 154.8 119.24 154.96 ;
      RECT 118.79 157.56 119.24 157.72 ;
      RECT 118.79 156.96 118.95 157.72 ;
      RECT 117.82 157.05 118.95 157.21 ;
      RECT 118.23 156.96 118.95 157.21 ;
      RECT 118.23 158.71 118.95 158.96 ;
      RECT 118.79 158.2 118.95 158.96 ;
      RECT 117.82 158.71 118.95 158.87 ;
      RECT 118.79 158.2 119.24 158.36 ;
      RECT 118.79 160.96 119.24 161.12 ;
      RECT 118.79 160.35 118.95 161.12 ;
      RECT 117.82 160.55 118.95 160.71 ;
      RECT 118.23 160.35 118.95 160.71 ;
      RECT 118.23 162.01 118.95 162.37 ;
      RECT 118.79 161.6 118.95 162.37 ;
      RECT 117.82 162.01 118.95 162.17 ;
      RECT 118.79 161.6 119.24 161.76 ;
      RECT 118.79 164.36 119.24 164.52 ;
      RECT 118.79 163.76 118.95 164.52 ;
      RECT 117.82 163.85 118.95 164.01 ;
      RECT 118.23 163.76 118.95 164.01 ;
      RECT 118.23 165.51 118.95 165.76 ;
      RECT 118.79 165 118.95 165.76 ;
      RECT 117.82 165.51 118.95 165.67 ;
      RECT 118.79 165 119.24 165.16 ;
      RECT 118.79 167.76 119.24 167.92 ;
      RECT 118.79 167.15 118.95 167.92 ;
      RECT 117.82 167.35 118.95 167.51 ;
      RECT 118.23 167.15 118.95 167.51 ;
      RECT 118.23 168.81 118.95 169.17 ;
      RECT 118.79 168.4 118.95 169.17 ;
      RECT 117.82 168.81 118.95 168.97 ;
      RECT 118.79 168.4 119.24 168.56 ;
      RECT 118.79 171.16 119.24 171.32 ;
      RECT 118.79 170.56 118.95 171.32 ;
      RECT 117.82 170.65 118.95 170.81 ;
      RECT 118.23 170.56 118.95 170.81 ;
      RECT 118.23 172.31 118.95 172.56 ;
      RECT 118.79 171.8 118.95 172.56 ;
      RECT 117.82 172.31 118.95 172.47 ;
      RECT 118.79 171.8 119.24 171.96 ;
      RECT 118.79 174.56 119.24 174.72 ;
      RECT 118.79 173.95 118.95 174.72 ;
      RECT 117.82 174.15 118.95 174.31 ;
      RECT 118.23 173.95 118.95 174.31 ;
      RECT 118.23 175.61 118.95 175.97 ;
      RECT 118.79 175.2 118.95 175.97 ;
      RECT 117.82 175.61 118.95 175.77 ;
      RECT 118.79 175.2 119.24 175.36 ;
      RECT 118.79 177.96 119.24 178.12 ;
      RECT 118.79 177.36 118.95 178.12 ;
      RECT 117.82 177.45 118.95 177.61 ;
      RECT 118.23 177.36 118.95 177.61 ;
      RECT 118.23 179.11 118.95 179.36 ;
      RECT 118.79 178.6 118.95 179.36 ;
      RECT 117.82 179.11 118.95 179.27 ;
      RECT 118.79 178.6 119.24 178.76 ;
      RECT 118.79 181.36 119.24 181.52 ;
      RECT 118.79 180.75 118.95 181.52 ;
      RECT 117.82 180.95 118.95 181.11 ;
      RECT 118.23 180.75 118.95 181.11 ;
      RECT 118.23 182.41 118.95 182.77 ;
      RECT 118.79 182 118.95 182.77 ;
      RECT 117.82 182.41 118.95 182.57 ;
      RECT 118.79 182 119.24 182.16 ;
      RECT 118.79 184.76 119.24 184.92 ;
      RECT 118.79 184.16 118.95 184.92 ;
      RECT 117.82 184.25 118.95 184.41 ;
      RECT 118.23 184.16 118.95 184.41 ;
      RECT 118.23 185.91 118.95 186.16 ;
      RECT 118.79 185.4 118.95 186.16 ;
      RECT 117.82 185.91 118.95 186.07 ;
      RECT 118.79 185.4 119.24 185.56 ;
      RECT 118.79 188.16 119.24 188.32 ;
      RECT 118.79 187.55 118.95 188.32 ;
      RECT 117.82 187.75 118.95 187.91 ;
      RECT 118.23 187.55 118.95 187.91 ;
      RECT 118.23 189.21 118.95 189.57 ;
      RECT 118.79 188.8 118.95 189.57 ;
      RECT 117.82 189.21 118.95 189.37 ;
      RECT 118.79 188.8 119.24 188.96 ;
      RECT 118.79 191.56 119.24 191.72 ;
      RECT 118.79 190.96 118.95 191.72 ;
      RECT 117.82 191.05 118.95 191.21 ;
      RECT 118.23 190.96 118.95 191.21 ;
      RECT 118.23 192.71 118.95 192.96 ;
      RECT 118.79 192.2 118.95 192.96 ;
      RECT 117.82 192.71 118.95 192.87 ;
      RECT 118.79 192.2 119.24 192.36 ;
      RECT 118.79 194.96 119.24 195.12 ;
      RECT 118.79 194.35 118.95 195.12 ;
      RECT 117.82 194.55 118.95 194.71 ;
      RECT 118.23 194.35 118.95 194.71 ;
      RECT 118.23 196.01 118.95 196.37 ;
      RECT 118.79 195.6 118.95 196.37 ;
      RECT 117.82 196.01 118.95 196.17 ;
      RECT 118.79 195.6 119.24 195.76 ;
      RECT 118.79 198.36 119.24 198.52 ;
      RECT 118.79 197.76 118.95 198.52 ;
      RECT 117.82 197.85 118.95 198.01 ;
      RECT 118.23 197.76 118.95 198.01 ;
      RECT 118.23 199.51 118.95 199.76 ;
      RECT 118.79 199 118.95 199.76 ;
      RECT 117.82 199.51 118.95 199.67 ;
      RECT 118.79 199 119.24 199.16 ;
      RECT 118.79 201.76 119.24 201.92 ;
      RECT 118.79 201.15 118.95 201.92 ;
      RECT 117.82 201.35 118.95 201.51 ;
      RECT 118.23 201.15 118.95 201.51 ;
      RECT 118.23 202.81 118.95 203.17 ;
      RECT 118.79 202.4 118.95 203.17 ;
      RECT 117.82 202.81 118.95 202.97 ;
      RECT 118.79 202.4 119.24 202.56 ;
      RECT 118.79 205.16 119.24 205.32 ;
      RECT 118.79 204.56 118.95 205.32 ;
      RECT 117.82 204.65 118.95 204.81 ;
      RECT 118.23 204.56 118.95 204.81 ;
      RECT 118.23 206.31 118.95 206.56 ;
      RECT 118.79 205.8 118.95 206.56 ;
      RECT 117.82 206.31 118.95 206.47 ;
      RECT 118.79 205.8 119.24 205.96 ;
      RECT 118.79 208.56 119.24 208.72 ;
      RECT 118.79 207.95 118.95 208.72 ;
      RECT 117.82 208.15 118.95 208.31 ;
      RECT 118.23 207.95 118.95 208.31 ;
      RECT 118.23 209.61 118.95 209.97 ;
      RECT 118.79 209.2 118.95 209.97 ;
      RECT 117.82 209.61 118.95 209.77 ;
      RECT 118.79 209.2 119.24 209.36 ;
      RECT 118.79 211.96 119.24 212.12 ;
      RECT 118.79 211.36 118.95 212.12 ;
      RECT 117.82 211.45 118.95 211.61 ;
      RECT 118.23 211.36 118.95 211.61 ;
      RECT 118.23 213.11 118.95 213.36 ;
      RECT 118.79 212.6 118.95 213.36 ;
      RECT 117.82 213.11 118.95 213.27 ;
      RECT 118.79 212.6 119.24 212.76 ;
      RECT 118.79 215.36 119.24 215.52 ;
      RECT 118.79 214.75 118.95 215.52 ;
      RECT 117.82 214.95 118.95 215.11 ;
      RECT 118.23 214.75 118.95 215.11 ;
      RECT 118.23 216.41 118.95 216.77 ;
      RECT 118.79 216 118.95 216.77 ;
      RECT 117.82 216.41 118.95 216.57 ;
      RECT 118.79 216 119.24 216.16 ;
      RECT 118.79 218.76 119.24 218.92 ;
      RECT 118.79 218.16 118.95 218.92 ;
      RECT 117.82 218.25 118.95 218.41 ;
      RECT 118.23 218.16 118.95 218.41 ;
      RECT 118.23 219.91 118.95 220.16 ;
      RECT 118.79 219.4 118.95 220.16 ;
      RECT 117.82 219.91 118.95 220.07 ;
      RECT 118.79 219.4 119.24 219.56 ;
      RECT 118.79 222.16 119.24 222.32 ;
      RECT 118.79 221.55 118.95 222.32 ;
      RECT 117.82 221.75 118.95 221.91 ;
      RECT 118.23 221.55 118.95 221.91 ;
      RECT 118.23 223.21 118.95 223.57 ;
      RECT 118.79 222.8 118.95 223.57 ;
      RECT 117.82 223.21 118.95 223.37 ;
      RECT 118.79 222.8 119.24 222.96 ;
      RECT 118.79 225.56 119.24 225.72 ;
      RECT 118.79 224.96 118.95 225.72 ;
      RECT 117.82 225.05 118.95 225.21 ;
      RECT 118.23 224.96 118.95 225.21 ;
      RECT 118.23 226.71 118.95 226.96 ;
      RECT 118.79 226.2 118.95 226.96 ;
      RECT 117.82 226.71 118.95 226.87 ;
      RECT 118.79 226.2 119.24 226.36 ;
      RECT 118.79 228.96 119.24 229.12 ;
      RECT 118.79 228.35 118.95 229.12 ;
      RECT 117.82 228.55 118.95 228.71 ;
      RECT 118.23 228.35 118.95 228.71 ;
      RECT 118.23 230.01 118.95 230.37 ;
      RECT 118.79 229.6 118.95 230.37 ;
      RECT 117.82 230.01 118.95 230.17 ;
      RECT 118.79 229.6 119.24 229.76 ;
      RECT 118.79 232.36 119.24 232.52 ;
      RECT 118.79 231.76 118.95 232.52 ;
      RECT 117.82 231.85 118.95 232.01 ;
      RECT 118.23 231.76 118.95 232.01 ;
      RECT 118.23 233.51 118.95 233.76 ;
      RECT 118.79 233 118.95 233.76 ;
      RECT 117.82 233.51 118.95 233.67 ;
      RECT 118.79 233 119.24 233.16 ;
      RECT 118.79 235.76 119.24 235.92 ;
      RECT 118.79 235.15 118.95 235.92 ;
      RECT 117.82 235.35 118.95 235.51 ;
      RECT 118.23 235.15 118.95 235.51 ;
      RECT 118.23 236.81 118.95 237.17 ;
      RECT 118.79 236.4 118.95 237.17 ;
      RECT 117.82 236.81 118.95 236.97 ;
      RECT 118.79 236.4 119.24 236.56 ;
      RECT 118.79 239.16 119.24 239.32 ;
      RECT 118.79 238.56 118.95 239.32 ;
      RECT 117.82 238.65 118.95 238.81 ;
      RECT 118.23 238.56 118.95 238.81 ;
      RECT 118.23 240.31 118.95 240.56 ;
      RECT 118.79 239.8 118.95 240.56 ;
      RECT 117.82 240.31 118.95 240.47 ;
      RECT 118.79 239.8 119.24 239.96 ;
      RECT 118.79 242.56 119.24 242.72 ;
      RECT 118.79 241.95 118.95 242.72 ;
      RECT 117.82 242.15 118.95 242.31 ;
      RECT 118.23 241.95 118.95 242.31 ;
      RECT 118.23 243.61 118.95 243.97 ;
      RECT 118.79 243.2 118.95 243.97 ;
      RECT 117.82 243.61 118.95 243.77 ;
      RECT 118.79 243.2 119.24 243.36 ;
      RECT 118.79 245.96 119.24 246.12 ;
      RECT 118.79 245.36 118.95 246.12 ;
      RECT 117.82 245.45 118.95 245.61 ;
      RECT 118.23 245.36 118.95 245.61 ;
      RECT 118.23 247.11 118.95 247.36 ;
      RECT 118.79 246.6 118.95 247.36 ;
      RECT 117.82 247.11 118.95 247.27 ;
      RECT 118.79 246.6 119.24 246.76 ;
      RECT 118.79 249.36 119.24 249.52 ;
      RECT 118.79 248.75 118.95 249.52 ;
      RECT 117.82 248.95 118.95 249.11 ;
      RECT 118.23 248.75 118.95 249.11 ;
      RECT 118.23 250.41 118.95 250.77 ;
      RECT 118.79 250 118.95 250.77 ;
      RECT 117.82 250.41 118.95 250.57 ;
      RECT 118.79 250 119.24 250.16 ;
      RECT 118.79 252.76 119.24 252.92 ;
      RECT 118.79 252.16 118.95 252.92 ;
      RECT 117.82 252.25 118.95 252.41 ;
      RECT 118.23 252.16 118.95 252.41 ;
      RECT 118.23 253.91 118.95 254.16 ;
      RECT 118.79 253.4 118.95 254.16 ;
      RECT 117.82 253.91 118.95 254.07 ;
      RECT 118.79 253.4 119.24 253.56 ;
      RECT 118.79 256.16 119.24 256.32 ;
      RECT 118.79 255.55 118.95 256.32 ;
      RECT 117.82 255.75 118.95 255.91 ;
      RECT 118.23 255.55 118.95 255.91 ;
      RECT 118.23 257.21 118.95 257.57 ;
      RECT 118.79 256.8 118.95 257.57 ;
      RECT 117.82 257.21 118.95 257.37 ;
      RECT 118.79 256.8 119.24 256.96 ;
      RECT 118.79 259.56 119.24 259.72 ;
      RECT 118.79 258.96 118.95 259.72 ;
      RECT 117.82 259.05 118.95 259.21 ;
      RECT 118.23 258.96 118.95 259.21 ;
      RECT 118.23 260.71 118.95 260.96 ;
      RECT 118.79 260.2 118.95 260.96 ;
      RECT 117.82 260.71 118.95 260.87 ;
      RECT 118.79 260.2 119.24 260.36 ;
      RECT 118.79 262.96 119.24 263.12 ;
      RECT 118.79 262.35 118.95 263.12 ;
      RECT 117.82 262.55 118.95 262.71 ;
      RECT 118.23 262.35 118.95 262.71 ;
      RECT 118.23 264.01 118.95 264.37 ;
      RECT 118.79 263.6 118.95 264.37 ;
      RECT 117.82 264.01 118.95 264.17 ;
      RECT 118.79 263.6 119.24 263.76 ;
      RECT 118.79 266.36 119.24 266.52 ;
      RECT 118.79 265.76 118.95 266.52 ;
      RECT 117.82 265.85 118.95 266.01 ;
      RECT 118.23 265.76 118.95 266.01 ;
      RECT 118.23 267.51 118.95 267.76 ;
      RECT 118.79 267 118.95 267.76 ;
      RECT 117.82 267.51 118.95 267.67 ;
      RECT 118.79 267 119.24 267.16 ;
      RECT 118.79 269.76 119.24 269.92 ;
      RECT 118.79 269.15 118.95 269.92 ;
      RECT 117.82 269.35 118.95 269.51 ;
      RECT 118.23 269.15 118.95 269.51 ;
      RECT 118.23 270.81 118.95 271.17 ;
      RECT 118.79 270.4 118.95 271.17 ;
      RECT 117.82 270.81 118.95 270.97 ;
      RECT 118.79 270.4 119.24 270.56 ;
      RECT 118.79 273.16 119.24 273.32 ;
      RECT 118.79 272.56 118.95 273.32 ;
      RECT 117.82 272.65 118.95 272.81 ;
      RECT 118.23 272.56 118.95 272.81 ;
      RECT 118.23 274.31 118.95 274.56 ;
      RECT 118.79 273.8 118.95 274.56 ;
      RECT 117.82 274.31 118.95 274.47 ;
      RECT 118.79 273.8 119.24 273.96 ;
      RECT 118.79 276.56 119.24 276.72 ;
      RECT 118.79 275.95 118.95 276.72 ;
      RECT 117.82 276.15 118.95 276.31 ;
      RECT 118.23 275.95 118.95 276.31 ;
      RECT 118.23 277.61 118.95 277.97 ;
      RECT 118.79 277.2 118.95 277.97 ;
      RECT 117.82 277.61 118.95 277.77 ;
      RECT 118.79 277.2 119.24 277.36 ;
      RECT 118.79 279.96 119.24 280.12 ;
      RECT 118.79 279.36 118.95 280.12 ;
      RECT 117.82 279.45 118.95 279.61 ;
      RECT 118.23 279.36 118.95 279.61 ;
      RECT 118.23 281.11 118.95 281.36 ;
      RECT 118.79 280.6 118.95 281.36 ;
      RECT 117.82 281.11 118.95 281.27 ;
      RECT 118.79 280.6 119.24 280.76 ;
      RECT 118.79 283.36 119.24 283.52 ;
      RECT 118.79 282.75 118.95 283.52 ;
      RECT 117.82 282.95 118.95 283.11 ;
      RECT 118.23 282.75 118.95 283.11 ;
      RECT 118.23 284.41 118.95 284.77 ;
      RECT 118.79 284 118.95 284.77 ;
      RECT 117.82 284.41 118.95 284.57 ;
      RECT 118.79 284 119.24 284.16 ;
      RECT 118.79 286.76 119.24 286.92 ;
      RECT 118.79 286.16 118.95 286.92 ;
      RECT 117.82 286.25 118.95 286.41 ;
      RECT 118.23 286.16 118.95 286.41 ;
      RECT 118.23 287.91 118.95 288.16 ;
      RECT 118.79 287.4 118.95 288.16 ;
      RECT 117.82 287.91 118.95 288.07 ;
      RECT 118.79 287.4 119.24 287.56 ;
      RECT 118.79 290.16 119.24 290.32 ;
      RECT 118.79 289.55 118.95 290.32 ;
      RECT 117.82 289.75 118.95 289.91 ;
      RECT 118.23 289.55 118.95 289.91 ;
      RECT 118.23 291.21 118.95 291.57 ;
      RECT 118.79 290.8 118.95 291.57 ;
      RECT 117.82 291.21 118.95 291.37 ;
      RECT 118.79 290.8 119.24 290.96 ;
      RECT 118.79 293.56 119.24 293.72 ;
      RECT 118.79 292.96 118.95 293.72 ;
      RECT 117.82 293.05 118.95 293.21 ;
      RECT 118.23 292.96 118.95 293.21 ;
      RECT 118.23 294.71 118.95 294.96 ;
      RECT 118.79 294.2 118.95 294.96 ;
      RECT 117.82 294.71 118.95 294.87 ;
      RECT 118.79 294.2 119.24 294.36 ;
      RECT 118.79 296.96 119.24 297.12 ;
      RECT 118.79 296.35 118.95 297.12 ;
      RECT 117.82 296.55 118.95 296.71 ;
      RECT 118.23 296.35 118.95 296.71 ;
      RECT 118.23 298.01 118.95 298.37 ;
      RECT 118.79 297.6 118.95 298.37 ;
      RECT 117.82 298.01 118.95 298.17 ;
      RECT 118.79 297.6 119.24 297.76 ;
      RECT 118.79 300.36 119.24 300.52 ;
      RECT 118.79 299.76 118.95 300.52 ;
      RECT 117.82 299.85 118.95 300.01 ;
      RECT 118.23 299.76 118.95 300.01 ;
      RECT 118.23 301.51 118.95 301.76 ;
      RECT 118.79 301 118.95 301.76 ;
      RECT 117.82 301.51 118.95 301.67 ;
      RECT 118.79 301 119.24 301.16 ;
      RECT 118.79 303.76 119.24 303.92 ;
      RECT 118.79 303.15 118.95 303.92 ;
      RECT 117.82 303.35 118.95 303.51 ;
      RECT 118.23 303.15 118.95 303.51 ;
      RECT 118.23 304.81 118.95 305.17 ;
      RECT 118.79 304.4 118.95 305.17 ;
      RECT 117.82 304.81 118.95 304.97 ;
      RECT 118.79 304.4 119.24 304.56 ;
      RECT 118.79 307.16 119.24 307.32 ;
      RECT 118.79 306.56 118.95 307.32 ;
      RECT 117.82 306.65 118.95 306.81 ;
      RECT 118.23 306.56 118.95 306.81 ;
      RECT 118.23 308.31 118.95 308.56 ;
      RECT 118.79 307.8 118.95 308.56 ;
      RECT 117.82 308.31 118.95 308.47 ;
      RECT 118.79 307.8 119.24 307.96 ;
      RECT 118.79 310.56 119.24 310.72 ;
      RECT 118.79 309.95 118.95 310.72 ;
      RECT 117.82 310.15 118.95 310.31 ;
      RECT 118.23 309.95 118.95 310.31 ;
      RECT 118.23 311.61 118.95 311.97 ;
      RECT 118.79 311.2 118.95 311.97 ;
      RECT 117.82 311.61 118.95 311.77 ;
      RECT 118.79 311.2 119.24 311.36 ;
      RECT 118.79 313.96 119.24 314.12 ;
      RECT 118.79 313.36 118.95 314.12 ;
      RECT 117.82 313.45 118.95 313.61 ;
      RECT 118.23 313.36 118.95 313.61 ;
      RECT 118.23 315.11 118.95 315.36 ;
      RECT 118.79 314.6 118.95 315.36 ;
      RECT 117.82 315.11 118.95 315.27 ;
      RECT 118.79 314.6 119.24 314.76 ;
      RECT 118.79 317.36 119.24 317.52 ;
      RECT 118.79 316.75 118.95 317.52 ;
      RECT 117.82 316.95 118.95 317.11 ;
      RECT 118.23 316.75 118.95 317.11 ;
      RECT 118.23 318.41 118.95 318.77 ;
      RECT 118.79 318 118.95 318.77 ;
      RECT 117.82 318.41 118.95 318.57 ;
      RECT 118.79 318 119.24 318.16 ;
      RECT 118.79 320.76 119.24 320.92 ;
      RECT 118.79 320.16 118.95 320.92 ;
      RECT 117.82 320.25 118.95 320.41 ;
      RECT 118.23 320.16 118.95 320.41 ;
      RECT 118.23 321.91 118.95 322.16 ;
      RECT 118.79 321.4 118.95 322.16 ;
      RECT 117.82 321.91 118.95 322.07 ;
      RECT 118.79 321.4 119.24 321.56 ;
      RECT 118.79 324.16 119.24 324.32 ;
      RECT 118.79 323.55 118.95 324.32 ;
      RECT 117.82 323.75 118.95 323.91 ;
      RECT 118.23 323.55 118.95 323.91 ;
      RECT 118.23 325.21 118.95 325.57 ;
      RECT 118.79 324.8 118.95 325.57 ;
      RECT 117.82 325.21 118.95 325.37 ;
      RECT 118.79 324.8 119.24 324.96 ;
      RECT 118.79 327.56 119.24 327.72 ;
      RECT 118.79 326.96 118.95 327.72 ;
      RECT 117.82 327.05 118.95 327.21 ;
      RECT 118.23 326.96 118.95 327.21 ;
      RECT 118.23 328.71 118.95 328.96 ;
      RECT 118.79 328.2 118.95 328.96 ;
      RECT 117.82 328.71 118.95 328.87 ;
      RECT 118.79 328.2 119.24 328.36 ;
      RECT 118.79 330.96 119.24 331.12 ;
      RECT 118.79 330.35 118.95 331.12 ;
      RECT 117.82 330.55 118.95 330.71 ;
      RECT 118.23 330.35 118.95 330.71 ;
      RECT 118.23 332.01 118.95 332.37 ;
      RECT 118.79 331.6 118.95 332.37 ;
      RECT 117.82 332.01 118.95 332.17 ;
      RECT 118.79 331.6 119.24 331.76 ;
      RECT 118.79 334.36 119.24 334.52 ;
      RECT 118.79 333.76 118.95 334.52 ;
      RECT 117.82 333.85 118.95 334.01 ;
      RECT 118.23 333.76 118.95 334.01 ;
      RECT 118.23 335.51 118.95 335.76 ;
      RECT 118.79 335 118.95 335.76 ;
      RECT 117.82 335.51 118.95 335.67 ;
      RECT 118.79 335 119.24 335.16 ;
      RECT 118.79 337.76 119.24 337.92 ;
      RECT 118.79 337.15 118.95 337.92 ;
      RECT 117.82 337.35 118.95 337.51 ;
      RECT 118.23 337.15 118.95 337.51 ;
      RECT 118.23 338.81 118.95 339.17 ;
      RECT 118.79 338.4 118.95 339.17 ;
      RECT 117.82 338.81 118.95 338.97 ;
      RECT 118.79 338.4 119.24 338.56 ;
      RECT 118.79 341.16 119.24 341.32 ;
      RECT 118.79 340.56 118.95 341.32 ;
      RECT 117.82 340.65 118.95 340.81 ;
      RECT 118.23 340.56 118.95 340.81 ;
      RECT 118.23 342.31 118.95 342.56 ;
      RECT 118.79 341.8 118.95 342.56 ;
      RECT 117.82 342.31 118.95 342.47 ;
      RECT 118.79 341.8 119.24 341.96 ;
      RECT 118.79 344.56 119.24 344.72 ;
      RECT 118.79 343.95 118.95 344.72 ;
      RECT 117.82 344.15 118.95 344.31 ;
      RECT 118.23 343.95 118.95 344.31 ;
      RECT 118.23 345.61 118.95 345.97 ;
      RECT 118.79 345.2 118.95 345.97 ;
      RECT 117.82 345.61 118.95 345.77 ;
      RECT 118.79 345.2 119.24 345.36 ;
      RECT 118.79 347.96 119.24 348.12 ;
      RECT 118.79 347.36 118.95 348.12 ;
      RECT 117.82 347.45 118.95 347.61 ;
      RECT 118.23 347.36 118.95 347.61 ;
      RECT 118.23 349.11 118.95 349.36 ;
      RECT 118.79 348.6 118.95 349.36 ;
      RECT 117.82 349.11 118.95 349.27 ;
      RECT 118.79 348.6 119.24 348.76 ;
      RECT 118.79 351.36 119.24 351.52 ;
      RECT 118.79 350.75 118.95 351.52 ;
      RECT 117.82 350.95 118.95 351.11 ;
      RECT 118.23 350.75 118.95 351.11 ;
      RECT 118.23 352.41 118.95 352.77 ;
      RECT 118.79 352 118.95 352.77 ;
      RECT 117.82 352.41 118.95 352.57 ;
      RECT 118.79 352 119.24 352.16 ;
      RECT 118.79 354.76 119.24 354.92 ;
      RECT 118.79 354.16 118.95 354.92 ;
      RECT 117.82 354.25 118.95 354.41 ;
      RECT 118.23 354.16 118.95 354.41 ;
      RECT 118.23 355.91 118.95 356.16 ;
      RECT 118.79 355.4 118.95 356.16 ;
      RECT 117.82 355.91 118.95 356.07 ;
      RECT 118.79 355.4 119.24 355.56 ;
      RECT 118.79 358.16 119.24 358.32 ;
      RECT 118.79 357.55 118.95 358.32 ;
      RECT 117.82 357.75 118.95 357.91 ;
      RECT 118.23 357.55 118.95 357.91 ;
      RECT 118.23 359.21 118.95 359.57 ;
      RECT 118.79 358.8 118.95 359.57 ;
      RECT 117.82 359.21 118.95 359.37 ;
      RECT 118.79 358.8 119.24 358.96 ;
      RECT 118.79 361.56 119.24 361.72 ;
      RECT 118.79 360.96 118.95 361.72 ;
      RECT 117.82 361.05 118.95 361.21 ;
      RECT 118.23 360.96 118.95 361.21 ;
      RECT 118.23 362.71 118.95 362.96 ;
      RECT 118.79 362.2 118.95 362.96 ;
      RECT 117.82 362.71 118.95 362.87 ;
      RECT 118.79 362.2 119.24 362.36 ;
      RECT 118.79 364.96 119.24 365.12 ;
      RECT 118.79 364.35 118.95 365.12 ;
      RECT 117.82 364.55 118.95 364.71 ;
      RECT 118.23 364.35 118.95 364.71 ;
      RECT 118.23 366.01 118.95 366.37 ;
      RECT 118.79 365.6 118.95 366.37 ;
      RECT 117.82 366.01 118.95 366.17 ;
      RECT 118.79 365.6 119.24 365.76 ;
      RECT 118.79 368.36 119.24 368.52 ;
      RECT 118.79 367.76 118.95 368.52 ;
      RECT 117.82 367.85 118.95 368.01 ;
      RECT 118.23 367.76 118.95 368.01 ;
      RECT 118.23 369.51 118.95 369.76 ;
      RECT 118.79 369 118.95 369.76 ;
      RECT 117.82 369.51 118.95 369.67 ;
      RECT 118.79 369 119.24 369.16 ;
      RECT 118.79 371.76 119.24 371.92 ;
      RECT 118.79 371.15 118.95 371.92 ;
      RECT 117.82 371.35 118.95 371.51 ;
      RECT 118.23 371.15 118.95 371.51 ;
      RECT 118.23 372.81 118.95 373.17 ;
      RECT 118.79 372.4 118.95 373.17 ;
      RECT 117.82 372.81 118.95 372.97 ;
      RECT 118.79 372.4 119.24 372.56 ;
      RECT 118.79 375.16 119.24 375.32 ;
      RECT 118.79 374.56 118.95 375.32 ;
      RECT 117.82 374.65 118.95 374.81 ;
      RECT 118.23 374.56 118.95 374.81 ;
      RECT 118.23 376.31 118.95 376.56 ;
      RECT 118.79 375.8 118.95 376.56 ;
      RECT 117.82 376.31 118.95 376.47 ;
      RECT 118.79 375.8 119.24 375.96 ;
      RECT 118.79 378.56 119.24 378.72 ;
      RECT 118.79 377.95 118.95 378.72 ;
      RECT 117.82 378.15 118.95 378.31 ;
      RECT 118.23 377.95 118.95 378.31 ;
      RECT 118.23 379.61 118.95 379.97 ;
      RECT 118.79 379.2 118.95 379.97 ;
      RECT 117.82 379.61 118.95 379.77 ;
      RECT 118.79 379.2 119.24 379.36 ;
      RECT 118.79 381.96 119.24 382.12 ;
      RECT 118.79 381.36 118.95 382.12 ;
      RECT 117.82 381.45 118.95 381.61 ;
      RECT 118.23 381.36 118.95 381.61 ;
      RECT 118.23 383.11 118.95 383.36 ;
      RECT 118.79 382.6 118.95 383.36 ;
      RECT 117.82 383.11 118.95 383.27 ;
      RECT 118.79 382.6 119.24 382.76 ;
      RECT 118.79 385.36 119.24 385.52 ;
      RECT 118.79 384.75 118.95 385.52 ;
      RECT 117.82 384.95 118.95 385.11 ;
      RECT 118.23 384.75 118.95 385.11 ;
      RECT 118.23 386.41 118.95 386.77 ;
      RECT 118.79 386 118.95 386.77 ;
      RECT 117.82 386.41 118.95 386.57 ;
      RECT 118.79 386 119.24 386.16 ;
      RECT 118.79 388.76 119.24 388.92 ;
      RECT 118.79 388.16 118.95 388.92 ;
      RECT 117.82 388.25 118.95 388.41 ;
      RECT 118.23 388.16 118.95 388.41 ;
      RECT 118.23 389.91 118.95 390.16 ;
      RECT 118.79 389.4 118.95 390.16 ;
      RECT 117.82 389.91 118.95 390.07 ;
      RECT 118.79 389.4 119.24 389.56 ;
      RECT 118.79 392.16 119.24 392.32 ;
      RECT 118.79 391.55 118.95 392.32 ;
      RECT 117.82 391.75 118.95 391.91 ;
      RECT 118.23 391.55 118.95 391.91 ;
      RECT 118.23 393.21 118.95 393.57 ;
      RECT 118.79 392.8 118.95 393.57 ;
      RECT 117.82 393.21 118.95 393.37 ;
      RECT 118.79 392.8 119.24 392.96 ;
      RECT 118.79 395.56 119.24 395.72 ;
      RECT 118.79 394.96 118.95 395.72 ;
      RECT 117.82 395.05 118.95 395.21 ;
      RECT 118.23 394.96 118.95 395.21 ;
      RECT 118.23 396.71 118.95 396.96 ;
      RECT 118.79 396.2 118.95 396.96 ;
      RECT 117.82 396.71 118.95 396.87 ;
      RECT 118.79 396.2 119.24 396.36 ;
      RECT 118.79 398.96 119.24 399.12 ;
      RECT 118.79 398.35 118.95 399.12 ;
      RECT 117.82 398.55 118.95 398.71 ;
      RECT 118.23 398.35 118.95 398.71 ;
      RECT 118.23 400.01 118.95 400.37 ;
      RECT 118.79 399.6 118.95 400.37 ;
      RECT 117.82 400.01 118.95 400.17 ;
      RECT 118.79 399.6 119.24 399.76 ;
      RECT 118.79 402.36 119.24 402.52 ;
      RECT 118.79 401.76 118.95 402.52 ;
      RECT 117.82 401.85 118.95 402.01 ;
      RECT 118.23 401.76 118.95 402.01 ;
      RECT 118.23 403.51 118.95 403.76 ;
      RECT 118.79 403 118.95 403.76 ;
      RECT 117.82 403.51 118.95 403.67 ;
      RECT 118.79 403 119.24 403.16 ;
      RECT 118.79 405.76 119.24 405.92 ;
      RECT 118.79 405.15 118.95 405.92 ;
      RECT 117.82 405.35 118.95 405.51 ;
      RECT 118.23 405.15 118.95 405.51 ;
      RECT 118.23 406.81 118.95 407.17 ;
      RECT 118.79 406.4 118.95 407.17 ;
      RECT 117.82 406.81 118.95 406.97 ;
      RECT 118.79 406.4 119.24 406.56 ;
      RECT 118.79 409.16 119.24 409.32 ;
      RECT 118.79 408.56 118.95 409.32 ;
      RECT 117.82 408.65 118.95 408.81 ;
      RECT 118.23 408.56 118.95 408.81 ;
      RECT 118.23 410.31 118.95 410.56 ;
      RECT 118.79 409.8 118.95 410.56 ;
      RECT 117.82 410.31 118.95 410.47 ;
      RECT 118.79 409.8 119.24 409.96 ;
      RECT 118.79 412.56 119.24 412.72 ;
      RECT 118.79 411.95 118.95 412.72 ;
      RECT 117.82 412.15 118.95 412.31 ;
      RECT 118.23 411.95 118.95 412.31 ;
      RECT 118.23 413.61 118.95 413.97 ;
      RECT 118.79 413.2 118.95 413.97 ;
      RECT 117.82 413.61 118.95 413.77 ;
      RECT 118.79 413.2 119.24 413.36 ;
      RECT 118.79 415.96 119.24 416.12 ;
      RECT 118.79 415.36 118.95 416.12 ;
      RECT 117.82 415.45 118.95 415.61 ;
      RECT 118.23 415.36 118.95 415.61 ;
      RECT 118.23 417.11 118.95 417.36 ;
      RECT 118.79 416.6 118.95 417.36 ;
      RECT 117.82 417.11 118.95 417.27 ;
      RECT 118.79 416.6 119.24 416.76 ;
      RECT 118.79 419.36 119.24 419.52 ;
      RECT 118.79 418.75 118.95 419.52 ;
      RECT 117.82 418.95 118.95 419.11 ;
      RECT 118.23 418.75 118.95 419.11 ;
      RECT 118.23 420.41 118.95 420.77 ;
      RECT 118.79 420 118.95 420.77 ;
      RECT 117.82 420.41 118.95 420.57 ;
      RECT 118.79 420 119.24 420.16 ;
      RECT 118.79 422.76 119.24 422.92 ;
      RECT 118.79 422.16 118.95 422.92 ;
      RECT 117.82 422.25 118.95 422.41 ;
      RECT 118.23 422.16 118.95 422.41 ;
      RECT 118.23 423.91 118.95 424.16 ;
      RECT 118.79 423.4 118.95 424.16 ;
      RECT 117.82 423.91 118.95 424.07 ;
      RECT 118.79 423.4 119.24 423.56 ;
      RECT 118.79 426.16 119.24 426.32 ;
      RECT 118.79 425.55 118.95 426.32 ;
      RECT 117.82 425.75 118.95 425.91 ;
      RECT 118.23 425.55 118.95 425.91 ;
      RECT 118.23 427.21 118.95 427.57 ;
      RECT 118.79 426.8 118.95 427.57 ;
      RECT 117.82 427.21 118.95 427.37 ;
      RECT 118.79 426.8 119.24 426.96 ;
      RECT 118.79 429.56 119.24 429.72 ;
      RECT 118.79 428.96 118.95 429.72 ;
      RECT 117.82 429.05 118.95 429.21 ;
      RECT 118.23 428.96 118.95 429.21 ;
      RECT 118.23 430.71 118.95 430.96 ;
      RECT 118.79 430.2 118.95 430.96 ;
      RECT 117.82 430.71 118.95 430.87 ;
      RECT 118.79 430.2 119.24 430.36 ;
      RECT 118.79 432.96 119.24 433.12 ;
      RECT 118.79 432.35 118.95 433.12 ;
      RECT 117.82 432.55 118.95 432.71 ;
      RECT 118.23 432.35 118.95 432.71 ;
      RECT 118.23 434.01 118.95 434.37 ;
      RECT 118.79 433.6 118.95 434.37 ;
      RECT 117.82 434.01 118.95 434.17 ;
      RECT 118.79 433.6 119.24 433.76 ;
      RECT 118.79 436.36 119.24 436.52 ;
      RECT 118.79 435.76 118.95 436.52 ;
      RECT 117.82 435.85 118.95 436.01 ;
      RECT 118.23 435.76 118.95 436.01 ;
      RECT 118.23 437.51 118.95 437.76 ;
      RECT 118.79 437 118.95 437.76 ;
      RECT 117.82 437.51 118.95 437.67 ;
      RECT 118.79 437 119.24 437.16 ;
      RECT 118.79 439.76 119.24 439.92 ;
      RECT 118.79 439.15 118.95 439.92 ;
      RECT 117.82 439.35 118.95 439.51 ;
      RECT 118.23 439.15 118.95 439.51 ;
      RECT 118.23 440.81 118.95 441.17 ;
      RECT 118.79 440.4 118.95 441.17 ;
      RECT 117.82 440.81 118.95 440.97 ;
      RECT 118.79 440.4 119.24 440.56 ;
      RECT 118.79 443.16 119.24 443.32 ;
      RECT 118.79 442.56 118.95 443.32 ;
      RECT 117.82 442.65 118.95 442.81 ;
      RECT 118.23 442.56 118.95 442.81 ;
      RECT 118.23 444.31 118.95 444.56 ;
      RECT 118.79 443.8 118.95 444.56 ;
      RECT 117.82 444.31 118.95 444.47 ;
      RECT 118.79 443.8 119.24 443.96 ;
      RECT 118.79 446.56 119.24 446.72 ;
      RECT 118.79 445.95 118.95 446.72 ;
      RECT 117.82 446.15 118.95 446.31 ;
      RECT 118.23 445.95 118.95 446.31 ;
      RECT 118.23 447.61 118.95 447.97 ;
      RECT 118.79 447.2 118.95 447.97 ;
      RECT 117.82 447.61 118.95 447.77 ;
      RECT 118.79 447.2 119.24 447.36 ;
      RECT 118.79 449.96 119.24 450.12 ;
      RECT 118.79 449.36 118.95 450.12 ;
      RECT 117.82 449.45 118.95 449.61 ;
      RECT 118.23 449.36 118.95 449.61 ;
      RECT 118.23 451.11 118.95 451.36 ;
      RECT 118.79 450.6 118.95 451.36 ;
      RECT 117.82 451.11 118.95 451.27 ;
      RECT 118.79 450.6 119.24 450.76 ;
      RECT 118.79 453.36 119.24 453.52 ;
      RECT 118.79 452.75 118.95 453.52 ;
      RECT 117.82 452.95 118.95 453.11 ;
      RECT 118.23 452.75 118.95 453.11 ;
      RECT 118.23 454.41 118.95 454.77 ;
      RECT 118.79 454 118.95 454.77 ;
      RECT 117.82 454.41 118.95 454.57 ;
      RECT 118.79 454 119.24 454.16 ;
      RECT 118.79 456.76 119.24 456.92 ;
      RECT 118.79 456.16 118.95 456.92 ;
      RECT 117.82 456.25 118.95 456.41 ;
      RECT 118.23 456.16 118.95 456.41 ;
      RECT 118.23 457.91 118.95 458.16 ;
      RECT 118.79 457.4 118.95 458.16 ;
      RECT 117.82 457.91 118.95 458.07 ;
      RECT 118.79 457.4 119.24 457.56 ;
      RECT 118.79 460.16 119.24 460.32 ;
      RECT 118.79 459.55 118.95 460.32 ;
      RECT 117.82 459.75 118.95 459.91 ;
      RECT 118.23 459.55 118.95 459.91 ;
      RECT 118.23 461.21 118.95 461.57 ;
      RECT 118.79 460.8 118.95 461.57 ;
      RECT 117.82 461.21 118.95 461.37 ;
      RECT 118.79 460.8 119.24 460.96 ;
      RECT 118.79 463.56 119.24 463.72 ;
      RECT 118.79 462.96 118.95 463.72 ;
      RECT 117.82 463.05 118.95 463.21 ;
      RECT 118.23 462.96 118.95 463.21 ;
      RECT 118.23 464.71 118.95 464.96 ;
      RECT 118.79 464.2 118.95 464.96 ;
      RECT 117.82 464.71 118.95 464.87 ;
      RECT 118.79 464.2 119.24 464.36 ;
      RECT 118.79 466.96 119.24 467.12 ;
      RECT 118.79 466.35 118.95 467.12 ;
      RECT 117.82 466.55 118.95 466.71 ;
      RECT 118.23 466.35 118.95 466.71 ;
      RECT 118.23 468.01 118.95 468.37 ;
      RECT 118.79 467.6 118.95 468.37 ;
      RECT 117.82 468.01 118.95 468.17 ;
      RECT 118.79 467.6 119.24 467.76 ;
      RECT 118.79 470.36 119.24 470.52 ;
      RECT 118.79 469.76 118.95 470.52 ;
      RECT 117.82 469.85 118.95 470.01 ;
      RECT 118.23 469.76 118.95 470.01 ;
      RECT 118.23 471.51 118.95 471.76 ;
      RECT 118.79 471 118.95 471.76 ;
      RECT 117.82 471.51 118.95 471.67 ;
      RECT 118.79 471 119.24 471.16 ;
      RECT 118.79 473.76 119.24 473.92 ;
      RECT 118.79 473.15 118.95 473.92 ;
      RECT 117.82 473.35 118.95 473.51 ;
      RECT 118.23 473.15 118.95 473.51 ;
      RECT 118.23 474.81 118.95 475.17 ;
      RECT 118.79 474.4 118.95 475.17 ;
      RECT 117.82 474.81 118.95 474.97 ;
      RECT 118.79 474.4 119.24 474.56 ;
      RECT 118.79 477.16 119.24 477.32 ;
      RECT 118.79 476.56 118.95 477.32 ;
      RECT 117.82 476.65 118.95 476.81 ;
      RECT 118.23 476.56 118.95 476.81 ;
      RECT 118.23 478.31 118.95 478.56 ;
      RECT 118.79 477.8 118.95 478.56 ;
      RECT 117.82 478.31 118.95 478.47 ;
      RECT 118.79 477.8 119.24 477.96 ;
      RECT 118.79 480.56 119.24 480.72 ;
      RECT 118.79 479.95 118.95 480.72 ;
      RECT 117.82 480.15 118.95 480.31 ;
      RECT 118.23 479.95 118.95 480.31 ;
      RECT 118.23 481.61 118.95 481.97 ;
      RECT 118.79 481.2 118.95 481.97 ;
      RECT 117.82 481.61 118.95 481.77 ;
      RECT 118.79 481.2 119.24 481.36 ;
      RECT 118.79 483.96 119.24 484.12 ;
      RECT 118.79 483.36 118.95 484.12 ;
      RECT 117.82 483.45 118.95 483.61 ;
      RECT 118.23 483.36 118.95 483.61 ;
      RECT 118.23 485.11 118.95 485.36 ;
      RECT 118.79 484.6 118.95 485.36 ;
      RECT 117.82 485.11 118.95 485.27 ;
      RECT 118.79 484.6 119.24 484.76 ;
      RECT 118.79 487.36 119.24 487.52 ;
      RECT 118.79 486.75 118.95 487.52 ;
      RECT 117.82 486.95 118.95 487.11 ;
      RECT 118.23 486.75 118.95 487.11 ;
      RECT 118.23 488.41 118.95 488.77 ;
      RECT 118.79 488 118.95 488.77 ;
      RECT 117.82 488.41 118.95 488.57 ;
      RECT 118.79 488 119.24 488.16 ;
      RECT 118.79 490.76 119.24 490.92 ;
      RECT 118.79 490.16 118.95 490.92 ;
      RECT 117.82 490.25 118.95 490.41 ;
      RECT 118.23 490.16 118.95 490.41 ;
      RECT 118.23 491.91 118.95 492.16 ;
      RECT 118.79 491.4 118.95 492.16 ;
      RECT 117.82 491.91 118.95 492.07 ;
      RECT 118.79 491.4 119.24 491.56 ;
      RECT 118.79 494.16 119.24 494.32 ;
      RECT 118.79 493.55 118.95 494.32 ;
      RECT 117.82 493.75 118.95 493.91 ;
      RECT 118.23 493.55 118.95 493.91 ;
      RECT 118.23 495.21 118.95 495.57 ;
      RECT 118.79 494.8 118.95 495.57 ;
      RECT 117.82 495.21 118.95 495.37 ;
      RECT 118.79 494.8 119.24 494.96 ;
      RECT 118.79 497.56 119.24 497.72 ;
      RECT 118.79 496.96 118.95 497.72 ;
      RECT 117.82 497.05 118.95 497.21 ;
      RECT 118.23 496.96 118.95 497.21 ;
      RECT 118.23 498.71 118.95 498.96 ;
      RECT 118.79 498.2 118.95 498.96 ;
      RECT 117.82 498.71 118.95 498.87 ;
      RECT 118.79 498.2 119.24 498.36 ;
      RECT 118.79 500.96 119.24 501.12 ;
      RECT 118.79 500.35 118.95 501.12 ;
      RECT 117.82 500.55 118.95 500.71 ;
      RECT 118.23 500.35 118.95 500.71 ;
      RECT 118.23 502.01 118.95 502.37 ;
      RECT 118.79 501.6 118.95 502.37 ;
      RECT 117.82 502.01 118.95 502.17 ;
      RECT 118.79 501.6 119.24 501.76 ;
      RECT 118.79 504.36 119.24 504.52 ;
      RECT 118.79 503.76 118.95 504.52 ;
      RECT 117.82 503.85 118.95 504.01 ;
      RECT 118.23 503.76 118.95 504.01 ;
      RECT 117.17 55.09 118.43 55.25 ;
      RECT 118.27 49.77 118.43 55.25 ;
      RECT 118.27 49.77 119.15 49.93 ;
      RECT 118.99 32.48 119.15 49.93 ;
      RECT 118.33 45.9 119.15 46.06 ;
      RECT 118.33 36.23 119.15 36.39 ;
      RECT 118.27 32.48 119.15 32.64 ;
      RECT 118.27 27.04 118.43 32.64 ;
      RECT 117.17 27.04 118.43 27.2 ;
      RECT 117.07 26.46 119.09 26.62 ;
      RECT 118.93 25.35 119.09 26.62 ;
      RECT 118.85 22.91 119.01 25.51 ;
      RECT 118.85 56.46 119.01 59.14 ;
      RECT 118.93 55.49 119.09 56.62 ;
      RECT 117.07 55.49 119.09 55.65 ;
      RECT 118.53 25.79 118.77 26.07 ;
      RECT 118.53 21.94 118.69 26.07 ;
      RECT 118.53 21.94 118.81 22.18 ;
      RECT 118.59 15.28 118.75 22.18 ;
      RECT 117.63 15.28 117.79 20.88 ;
      RECT 116.67 15.28 116.83 20.88 ;
      RECT 116.67 17.14 118.75 17.3 ;
      RECT 118.59 59.87 118.75 66.77 ;
      RECT 117.63 61.17 117.79 66.77 ;
      RECT 116.67 61.17 116.83 66.77 ;
      RECT 116.67 64.75 118.75 64.91 ;
      RECT 118.53 59.87 118.81 60.11 ;
      RECT 118.53 56.02 118.69 60.11 ;
      RECT 118.53 56.02 118.77 56.3 ;
      RECT 116.67 35.91 118.75 36.07 ;
      RECT 118.59 32.85 118.75 36.07 ;
      RECT 117.63 27.43 117.79 36.07 ;
      RECT 116.67 32.85 116.83 36.07 ;
      RECT 116.73 27.43 117.79 27.59 ;
      RECT 116.73 23.41 116.89 27.59 ;
      RECT 116.73 26.14 117.89 26.3 ;
      RECT 117.73 25.01 117.89 26.3 ;
      RECT 116.73 25 116.93 26.3 ;
      RECT 117.73 21.38 117.89 23.81 ;
      RECT 116.77 21.38 116.93 23.55 ;
      RECT 116.77 21.38 117.89 21.54 ;
      RECT 116.77 60.51 117.89 60.67 ;
      RECT 117.73 58.24 117.89 60.67 ;
      RECT 116.77 58.5 116.93 60.67 ;
      RECT 116.73 55.81 116.89 58.64 ;
      RECT 117.73 55.81 117.89 57.09 ;
      RECT 116.71 55.81 116.93 57.09 ;
      RECT 116.71 55.81 117.89 55.97 ;
      RECT 116.71 54.64 116.87 57.09 ;
      RECT 116.71 54.64 117.79 54.8 ;
      RECT 117.63 46.22 117.79 54.8 ;
      RECT 118.59 46.22 118.75 49.44 ;
      RECT 116.67 46.22 116.83 49.44 ;
      RECT 116.67 46.22 118.75 46.38 ;
      RECT 118.03 12.8 118.69 13.06 ;
      RECT 118.45 12.19 118.69 13.06 ;
      RECT 118.51 41.08 118.67 45.17 ;
      RECT 118.35 41.08 118.67 41.24 ;
      RECT 118.21 21.06 118.37 26.28 ;
      RECT 117.25 24.37 117.41 25.98 ;
      RECT 117.05 24.37 118.37 24.53 ;
      RECT 117.05 23.67 117.21 24.53 ;
      RECT 117.05 23.67 117.41 23.83 ;
      RECT 117.25 21.7 117.41 23.83 ;
      RECT 116.55 21.06 118.43 21.22 ;
      RECT 116.55 60.83 118.43 60.99 ;
      RECT 118.21 55.81 118.37 60.99 ;
      RECT 117.25 58.22 117.41 60.35 ;
      RECT 117.05 58.22 117.41 58.38 ;
      RECT 117.05 57.25 117.21 58.38 ;
      RECT 117.05 57.25 118.37 57.41 ;
      RECT 117.25 56.13 117.41 57.41 ;
      RECT 118.11 14.52 118.27 16.86 ;
      RECT 118.24 13.22 118.4 14.84 ;
      RECT 118.11 32.85 118.27 35.75 ;
      RECT 117.95 31.09 118.11 33.01 ;
      RECT 117.95 49.44 118.11 51.3 ;
      RECT 118.11 46.54 118.27 49.6 ;
      RECT 118.03 38.57 118.19 45.17 ;
      RECT 117.73 38.57 118.19 38.73 ;
      RECT 117.73 36.23 117.89 38.73 ;
      RECT 117.37 36.23 118.05 36.39 ;
      RECT 117.25 45.9 118.05 46.06 ;
      RECT 117.25 44.89 117.41 46.06 ;
      RECT 117.23 38.57 117.39 45.17 ;
      RECT 117.63 10.09 117.79 14.2 ;
      RECT 116.73 12.9 117.79 13.06 ;
      RECT 116.73 12.19 116.89 13.06 ;
      RECT 117.15 14.52 117.31 16.86 ;
      RECT 117.02 13.22 117.18 14.84 ;
      RECT 117.15 31.09 117.31 35.75 ;
      RECT 117.05 32.25 117.31 32.53 ;
      RECT 117.11 49.75 117.31 51.3 ;
      RECT 117.15 46.54 117.31 51.3 ;
      RECT 116.71 49.6 116.87 51.7 ;
      RECT 116.27 49.6 116.87 49.76 ;
      RECT 116.27 32.06 116.43 49.76 ;
      RECT 116.27 45.9 117.09 46.06 ;
      RECT 116.27 36.23 117.09 36.39 ;
      RECT 116.27 32.06 116.87 32.22 ;
      RECT 116.71 30.54 116.87 32.22 ;
      RECT 116.75 41.08 116.91 45.17 ;
      RECT 116.75 41.08 117.07 41.24 ;
      RECT 115.84 504.68 116.76 504.84 ;
      RECT 106.83 493.56 107.39 504.76 ;
      RECT 116.25 69.48 116.41 504.84 ;
      RECT 105.98 503.63 109.21 504.59 ;
      RECT 105.98 503.8 115.11 504.36 ;
      RECT 105.97 504.03 116.41 504.19 ;
      RECT 110.57 501.5 113.2 504.36 ;
      RECT 116.25 502.93 116.76 503.09 ;
      RECT 115.35 501.91 115.51 502.69 ;
      RECT 105.98 501.53 109.06 502.49 ;
      RECT 110.57 501.91 116.41 502.07 ;
      RECT 110.57 501.59 116.41 501.75 ;
      RECT 116.25 501.28 116.76 501.44 ;
      RECT 110.57 498.36 113.2 501.22 ;
      RECT 105.98 500.23 109.06 501.19 ;
      RECT 110.57 500.97 116.41 501.13 ;
      RECT 110.57 500.65 116.41 500.81 ;
      RECT 115.35 500.03 115.51 500.81 ;
      RECT 105.98 498.13 109.21 499.09 ;
      RECT 105.98 498.36 115.11 498.92 ;
      RECT 105.97 498.53 116.41 498.69 ;
      RECT 115.84 497.88 116.41 498.04 ;
      RECT 105.98 496.83 109.21 497.79 ;
      RECT 105.98 497 115.11 497.56 ;
      RECT 105.97 497.23 116.41 497.39 ;
      RECT 110.57 494.7 113.2 497.56 ;
      RECT 115.35 495.11 115.51 495.89 ;
      RECT 105.98 494.73 109.06 495.69 ;
      RECT 110.57 495.11 116.41 495.27 ;
      RECT 110.57 494.79 116.41 494.95 ;
      RECT 110.57 491.56 113.2 494.42 ;
      RECT 110.57 494.17 116.41 494.33 ;
      RECT 102.82 493.42 103.1 494.16 ;
      RECT 106.83 493.56 108.71 494.12 ;
      RECT 105.37 493.56 108.71 494.11 ;
      RECT 103.49 493.46 105.37 494.02 ;
      RECT 110.57 493.85 116.41 494.01 ;
      RECT 115.35 493.23 115.51 494.01 ;
      RECT 102.82 493.47 105.37 494.02 ;
      RECT 109.21 491.56 115.11 492.12 ;
      RECT 109.21 491.73 116.41 491.89 ;
      RECT 115.84 491.08 116.41 491.24 ;
      RECT 106.83 479.96 107.39 491.16 ;
      RECT 105.98 490.03 109.21 490.99 ;
      RECT 105.98 490.2 115.11 490.76 ;
      RECT 105.97 490.43 116.41 490.59 ;
      RECT 110.57 487.9 113.2 490.76 ;
      RECT 115.35 488.31 115.51 489.09 ;
      RECT 105.98 487.93 109.06 488.89 ;
      RECT 110.57 488.31 116.41 488.47 ;
      RECT 110.57 487.99 116.41 488.15 ;
      RECT 110.57 484.76 113.2 487.62 ;
      RECT 105.98 486.63 109.06 487.59 ;
      RECT 110.57 487.37 116.41 487.53 ;
      RECT 110.57 487.05 116.41 487.21 ;
      RECT 115.35 486.43 115.51 487.21 ;
      RECT 105.98 484.53 109.21 485.49 ;
      RECT 105.98 484.76 115.11 485.32 ;
      RECT 105.97 484.93 116.41 485.09 ;
      RECT 115.84 484.28 116.41 484.44 ;
      RECT 105.98 483.23 109.21 484.19 ;
      RECT 105.98 483.4 115.11 483.96 ;
      RECT 105.97 483.63 116.41 483.79 ;
      RECT 110.57 481.1 113.2 483.96 ;
      RECT 115.35 481.51 115.51 482.29 ;
      RECT 105.98 481.13 109.06 482.09 ;
      RECT 110.57 481.51 116.41 481.67 ;
      RECT 110.57 481.19 116.41 481.35 ;
      RECT 110.57 477.96 113.2 480.82 ;
      RECT 110.57 480.57 116.41 480.73 ;
      RECT 102.82 479.82 103.1 480.56 ;
      RECT 106.83 479.96 108.71 480.52 ;
      RECT 105.37 479.96 108.71 480.51 ;
      RECT 103.49 479.86 105.37 480.42 ;
      RECT 110.57 480.25 116.41 480.41 ;
      RECT 115.35 479.63 115.51 480.41 ;
      RECT 102.82 479.87 105.37 480.42 ;
      RECT 109.21 477.96 115.11 478.52 ;
      RECT 109.21 478.13 116.41 478.29 ;
      RECT 115.84 477.48 116.41 477.64 ;
      RECT 106.83 466.36 107.39 477.56 ;
      RECT 105.98 476.43 109.21 477.39 ;
      RECT 105.98 476.6 115.11 477.16 ;
      RECT 105.97 476.83 116.41 476.99 ;
      RECT 110.57 474.3 113.2 477.16 ;
      RECT 115.35 474.71 115.51 475.49 ;
      RECT 105.98 474.33 109.06 475.29 ;
      RECT 110.57 474.71 116.41 474.87 ;
      RECT 110.57 474.39 116.41 474.55 ;
      RECT 110.57 471.16 113.2 474.02 ;
      RECT 105.98 473.03 109.06 473.99 ;
      RECT 110.57 473.77 116.41 473.93 ;
      RECT 110.57 473.45 116.41 473.61 ;
      RECT 115.35 472.83 115.51 473.61 ;
      RECT 105.98 470.93 109.21 471.89 ;
      RECT 105.98 471.16 115.11 471.72 ;
      RECT 105.97 471.33 116.41 471.49 ;
      RECT 115.84 470.68 116.41 470.84 ;
      RECT 105.98 469.63 109.21 470.59 ;
      RECT 105.98 469.8 115.11 470.36 ;
      RECT 105.97 470.03 116.41 470.19 ;
      RECT 110.57 467.5 113.2 470.36 ;
      RECT 115.35 467.91 115.51 468.69 ;
      RECT 105.98 467.53 109.06 468.49 ;
      RECT 110.57 467.91 116.41 468.07 ;
      RECT 110.57 467.59 116.41 467.75 ;
      RECT 110.57 464.36 113.2 467.22 ;
      RECT 110.57 466.97 116.41 467.13 ;
      RECT 102.82 466.22 103.1 466.96 ;
      RECT 106.83 466.36 108.71 466.92 ;
      RECT 105.37 466.36 108.71 466.91 ;
      RECT 103.49 466.26 105.37 466.82 ;
      RECT 110.57 466.65 116.41 466.81 ;
      RECT 115.35 466.03 115.51 466.81 ;
      RECT 102.82 466.27 105.37 466.82 ;
      RECT 109.21 464.36 115.11 464.92 ;
      RECT 109.21 464.53 116.41 464.69 ;
      RECT 115.84 463.88 116.41 464.04 ;
      RECT 106.83 452.76 107.39 463.96 ;
      RECT 105.98 462.83 109.21 463.79 ;
      RECT 105.98 463 115.11 463.56 ;
      RECT 105.97 463.23 116.41 463.39 ;
      RECT 110.57 460.7 113.2 463.56 ;
      RECT 115.35 461.11 115.51 461.89 ;
      RECT 105.98 460.73 109.06 461.69 ;
      RECT 110.57 461.11 116.41 461.27 ;
      RECT 110.57 460.79 116.41 460.95 ;
      RECT 110.57 457.56 113.2 460.42 ;
      RECT 105.98 459.43 109.06 460.39 ;
      RECT 110.57 460.17 116.41 460.33 ;
      RECT 110.57 459.85 116.41 460.01 ;
      RECT 115.35 459.23 115.51 460.01 ;
      RECT 105.98 457.33 109.21 458.29 ;
      RECT 105.98 457.56 115.11 458.12 ;
      RECT 105.97 457.73 116.41 457.89 ;
      RECT 115.84 457.08 116.41 457.24 ;
      RECT 105.98 456.03 109.21 456.99 ;
      RECT 105.98 456.2 115.11 456.76 ;
      RECT 105.97 456.43 116.41 456.59 ;
      RECT 110.57 453.9 113.2 456.76 ;
      RECT 115.35 454.31 115.51 455.09 ;
      RECT 105.98 453.93 109.06 454.89 ;
      RECT 110.57 454.31 116.41 454.47 ;
      RECT 110.57 453.99 116.41 454.15 ;
      RECT 110.57 450.76 113.2 453.62 ;
      RECT 110.57 453.37 116.41 453.53 ;
      RECT 102.82 452.62 103.1 453.36 ;
      RECT 106.83 452.76 108.71 453.32 ;
      RECT 105.37 452.76 108.71 453.31 ;
      RECT 103.49 452.66 105.37 453.22 ;
      RECT 110.57 453.05 116.41 453.21 ;
      RECT 115.35 452.43 115.51 453.21 ;
      RECT 102.82 452.67 105.37 453.22 ;
      RECT 109.21 450.76 115.11 451.32 ;
      RECT 109.21 450.93 116.41 451.09 ;
      RECT 115.84 450.28 116.41 450.44 ;
      RECT 106.83 439.16 107.39 450.36 ;
      RECT 105.98 449.23 109.21 450.19 ;
      RECT 105.98 449.4 115.11 449.96 ;
      RECT 105.97 449.63 116.41 449.79 ;
      RECT 110.57 447.1 113.2 449.96 ;
      RECT 115.35 447.51 115.51 448.29 ;
      RECT 105.98 447.13 109.06 448.09 ;
      RECT 110.57 447.51 116.41 447.67 ;
      RECT 110.57 447.19 116.41 447.35 ;
      RECT 110.57 443.96 113.2 446.82 ;
      RECT 105.98 445.83 109.06 446.79 ;
      RECT 110.57 446.57 116.41 446.73 ;
      RECT 110.57 446.25 116.41 446.41 ;
      RECT 115.35 445.63 115.51 446.41 ;
      RECT 105.98 443.73 109.21 444.69 ;
      RECT 105.98 443.96 115.11 444.52 ;
      RECT 105.97 444.13 116.41 444.29 ;
      RECT 115.84 443.48 116.41 443.64 ;
      RECT 105.98 442.43 109.21 443.39 ;
      RECT 105.98 442.6 115.11 443.16 ;
      RECT 105.97 442.83 116.41 442.99 ;
      RECT 110.57 440.3 113.2 443.16 ;
      RECT 115.35 440.71 115.51 441.49 ;
      RECT 105.98 440.33 109.06 441.29 ;
      RECT 110.57 440.71 116.41 440.87 ;
      RECT 110.57 440.39 116.41 440.55 ;
      RECT 110.57 437.16 113.2 440.02 ;
      RECT 110.57 439.77 116.41 439.93 ;
      RECT 102.82 439.02 103.1 439.76 ;
      RECT 106.83 439.16 108.71 439.72 ;
      RECT 105.37 439.16 108.71 439.71 ;
      RECT 103.49 439.06 105.37 439.62 ;
      RECT 110.57 439.45 116.41 439.61 ;
      RECT 115.35 438.83 115.51 439.61 ;
      RECT 102.82 439.07 105.37 439.62 ;
      RECT 109.21 437.16 115.11 437.72 ;
      RECT 109.21 437.33 116.41 437.49 ;
      RECT 115.84 436.68 116.41 436.84 ;
      RECT 106.83 425.56 107.39 436.76 ;
      RECT 105.98 435.63 109.21 436.59 ;
      RECT 105.98 435.8 115.11 436.36 ;
      RECT 105.97 436.03 116.41 436.19 ;
      RECT 110.57 433.5 113.2 436.36 ;
      RECT 115.35 433.91 115.51 434.69 ;
      RECT 105.98 433.53 109.06 434.49 ;
      RECT 110.57 433.91 116.41 434.07 ;
      RECT 110.57 433.59 116.41 433.75 ;
      RECT 110.57 430.36 113.2 433.22 ;
      RECT 105.98 432.23 109.06 433.19 ;
      RECT 110.57 432.97 116.41 433.13 ;
      RECT 110.57 432.65 116.41 432.81 ;
      RECT 115.35 432.03 115.51 432.81 ;
      RECT 105.98 430.13 109.21 431.09 ;
      RECT 105.98 430.36 115.11 430.92 ;
      RECT 105.97 430.53 116.41 430.69 ;
      RECT 115.84 429.88 116.41 430.04 ;
      RECT 105.98 428.83 109.21 429.79 ;
      RECT 105.98 429 115.11 429.56 ;
      RECT 105.97 429.23 116.41 429.39 ;
      RECT 110.57 426.7 113.2 429.56 ;
      RECT 115.35 427.11 115.51 427.89 ;
      RECT 105.98 426.73 109.06 427.69 ;
      RECT 110.57 427.11 116.41 427.27 ;
      RECT 110.57 426.79 116.41 426.95 ;
      RECT 110.57 423.56 113.2 426.42 ;
      RECT 110.57 426.17 116.41 426.33 ;
      RECT 102.82 425.42 103.1 426.16 ;
      RECT 106.83 425.56 108.71 426.12 ;
      RECT 105.37 425.56 108.71 426.11 ;
      RECT 103.49 425.46 105.37 426.02 ;
      RECT 110.57 425.85 116.41 426.01 ;
      RECT 115.35 425.23 115.51 426.01 ;
      RECT 102.82 425.47 105.37 426.02 ;
      RECT 109.21 423.56 115.11 424.12 ;
      RECT 109.21 423.73 116.41 423.89 ;
      RECT 115.84 423.08 116.41 423.24 ;
      RECT 106.83 411.96 107.39 423.16 ;
      RECT 105.98 422.03 109.21 422.99 ;
      RECT 105.98 422.2 115.11 422.76 ;
      RECT 105.97 422.43 116.41 422.59 ;
      RECT 110.57 419.9 113.2 422.76 ;
      RECT 115.35 420.31 115.51 421.09 ;
      RECT 105.98 419.93 109.06 420.89 ;
      RECT 110.57 420.31 116.41 420.47 ;
      RECT 110.57 419.99 116.41 420.15 ;
      RECT 110.57 416.76 113.2 419.62 ;
      RECT 105.98 418.63 109.06 419.59 ;
      RECT 110.57 419.37 116.41 419.53 ;
      RECT 110.57 419.05 116.41 419.21 ;
      RECT 115.35 418.43 115.51 419.21 ;
      RECT 105.98 416.53 109.21 417.49 ;
      RECT 105.98 416.76 115.11 417.32 ;
      RECT 105.97 416.93 116.41 417.09 ;
      RECT 115.84 416.28 116.41 416.44 ;
      RECT 105.98 415.23 109.21 416.19 ;
      RECT 105.98 415.4 115.11 415.96 ;
      RECT 105.97 415.63 116.41 415.79 ;
      RECT 110.57 413.1 113.2 415.96 ;
      RECT 115.35 413.51 115.51 414.29 ;
      RECT 105.98 413.13 109.06 414.09 ;
      RECT 110.57 413.51 116.41 413.67 ;
      RECT 110.57 413.19 116.41 413.35 ;
      RECT 110.57 409.96 113.2 412.82 ;
      RECT 110.57 412.57 116.41 412.73 ;
      RECT 102.82 411.82 103.1 412.56 ;
      RECT 106.83 411.96 108.71 412.52 ;
      RECT 105.37 411.96 108.71 412.51 ;
      RECT 103.49 411.86 105.37 412.42 ;
      RECT 110.57 412.25 116.41 412.41 ;
      RECT 115.35 411.63 115.51 412.41 ;
      RECT 102.82 411.87 105.37 412.42 ;
      RECT 109.21 409.96 115.11 410.52 ;
      RECT 109.21 410.13 116.41 410.29 ;
      RECT 115.84 409.48 116.41 409.64 ;
      RECT 106.83 398.36 107.39 409.56 ;
      RECT 105.98 408.43 109.21 409.39 ;
      RECT 105.98 408.6 115.11 409.16 ;
      RECT 105.97 408.83 116.41 408.99 ;
      RECT 110.57 406.3 113.2 409.16 ;
      RECT 115.35 406.71 115.51 407.49 ;
      RECT 105.98 406.33 109.06 407.29 ;
      RECT 110.57 406.71 116.41 406.87 ;
      RECT 110.57 406.39 116.41 406.55 ;
      RECT 110.57 403.16 113.2 406.02 ;
      RECT 105.98 405.03 109.06 405.99 ;
      RECT 110.57 405.77 116.41 405.93 ;
      RECT 110.57 405.45 116.41 405.61 ;
      RECT 115.35 404.83 115.51 405.61 ;
      RECT 105.98 402.93 109.21 403.89 ;
      RECT 105.98 403.16 115.11 403.72 ;
      RECT 105.97 403.33 116.41 403.49 ;
      RECT 115.84 402.68 116.41 402.84 ;
      RECT 105.98 401.63 109.21 402.59 ;
      RECT 105.98 401.8 115.11 402.36 ;
      RECT 105.97 402.03 116.41 402.19 ;
      RECT 110.57 399.5 113.2 402.36 ;
      RECT 115.35 399.91 115.51 400.69 ;
      RECT 105.98 399.53 109.06 400.49 ;
      RECT 110.57 399.91 116.41 400.07 ;
      RECT 110.57 399.59 116.41 399.75 ;
      RECT 110.57 396.36 113.2 399.22 ;
      RECT 110.57 398.97 116.41 399.13 ;
      RECT 102.82 398.22 103.1 398.96 ;
      RECT 105.37 398.36 108.71 398.92 ;
      RECT 103.49 398.26 105.37 398.82 ;
      RECT 110.57 398.65 116.41 398.81 ;
      RECT 115.35 398.03 115.51 398.81 ;
      RECT 102.82 398.27 105.37 398.82 ;
      RECT 109.21 396.36 115.11 396.92 ;
      RECT 109.21 396.53 116.41 396.69 ;
      RECT 115.84 395.88 116.41 396.04 ;
      RECT 106.83 384.76 107.39 395.96 ;
      RECT 105.98 394.83 109.21 395.79 ;
      RECT 105.98 395 115.11 395.56 ;
      RECT 105.97 395.23 116.41 395.39 ;
      RECT 110.57 392.7 113.2 395.56 ;
      RECT 115.35 393.11 115.51 393.89 ;
      RECT 105.98 392.73 109.06 393.69 ;
      RECT 110.57 393.11 116.41 393.27 ;
      RECT 110.57 392.79 116.41 392.95 ;
      RECT 110.57 389.56 113.2 392.42 ;
      RECT 105.98 391.43 109.06 392.39 ;
      RECT 110.57 392.17 116.41 392.33 ;
      RECT 110.57 391.85 116.41 392.01 ;
      RECT 115.35 391.23 115.51 392.01 ;
      RECT 105.98 389.33 109.21 390.29 ;
      RECT 105.98 389.56 115.11 390.12 ;
      RECT 105.97 389.73 116.41 389.89 ;
      RECT 115.84 389.08 116.41 389.24 ;
      RECT 105.98 388.03 109.21 388.99 ;
      RECT 105.98 388.2 115.11 388.76 ;
      RECT 105.97 388.43 116.41 388.59 ;
      RECT 110.57 385.9 113.2 388.76 ;
      RECT 115.35 386.31 115.51 387.09 ;
      RECT 105.98 385.93 109.06 386.89 ;
      RECT 110.57 386.31 116.41 386.47 ;
      RECT 110.57 385.99 116.41 386.15 ;
      RECT 110.57 382.76 113.2 385.62 ;
      RECT 110.57 385.37 116.41 385.53 ;
      RECT 102.82 384.62 103.1 385.36 ;
      RECT 106.83 384.76 108.71 385.32 ;
      RECT 105.37 384.76 108.71 385.31 ;
      RECT 103.49 384.66 105.37 385.22 ;
      RECT 110.57 385.05 116.41 385.21 ;
      RECT 115.35 384.43 115.51 385.21 ;
      RECT 102.82 384.67 105.37 385.22 ;
      RECT 109.21 382.76 115.11 383.32 ;
      RECT 109.21 382.93 116.41 383.09 ;
      RECT 115.84 382.28 116.41 382.44 ;
      RECT 106.83 371.16 107.39 382.36 ;
      RECT 105.98 381.23 109.21 382.19 ;
      RECT 105.98 381.4 115.11 381.96 ;
      RECT 105.97 381.63 116.41 381.79 ;
      RECT 110.57 379.1 113.2 381.96 ;
      RECT 115.35 379.51 115.51 380.29 ;
      RECT 105.98 379.13 109.06 380.09 ;
      RECT 110.57 379.51 116.41 379.67 ;
      RECT 110.57 379.19 116.41 379.35 ;
      RECT 110.57 375.96 113.2 378.82 ;
      RECT 105.98 377.83 109.06 378.79 ;
      RECT 110.57 378.57 116.41 378.73 ;
      RECT 110.57 378.25 116.41 378.41 ;
      RECT 115.35 377.63 115.51 378.41 ;
      RECT 105.98 375.73 109.21 376.69 ;
      RECT 105.98 375.96 115.11 376.52 ;
      RECT 105.97 376.13 116.41 376.29 ;
      RECT 115.84 375.48 116.41 375.64 ;
      RECT 105.98 374.43 109.21 375.39 ;
      RECT 105.98 374.6 115.11 375.16 ;
      RECT 105.97 374.83 116.41 374.99 ;
      RECT 110.57 372.3 113.2 375.16 ;
      RECT 115.35 372.71 115.51 373.49 ;
      RECT 105.98 372.33 109.06 373.29 ;
      RECT 110.57 372.71 116.41 372.87 ;
      RECT 110.57 372.39 116.41 372.55 ;
      RECT 110.57 369.16 113.2 372.02 ;
      RECT 110.57 371.77 116.41 371.93 ;
      RECT 102.82 371.02 103.1 371.76 ;
      RECT 106.83 371.16 108.71 371.72 ;
      RECT 105.37 371.16 108.71 371.71 ;
      RECT 103.49 371.06 105.37 371.62 ;
      RECT 110.57 371.45 116.41 371.61 ;
      RECT 115.35 370.83 115.51 371.61 ;
      RECT 102.82 371.07 105.37 371.62 ;
      RECT 109.21 369.16 115.11 369.72 ;
      RECT 109.21 369.33 116.41 369.49 ;
      RECT 115.84 368.68 116.41 368.84 ;
      RECT 106.83 357.56 107.39 368.76 ;
      RECT 105.98 367.63 109.21 368.59 ;
      RECT 105.98 367.8 115.11 368.36 ;
      RECT 105.97 368.03 116.41 368.19 ;
      RECT 110.57 365.5 113.2 368.36 ;
      RECT 115.35 365.91 115.51 366.69 ;
      RECT 105.98 365.53 109.06 366.49 ;
      RECT 110.57 365.91 116.41 366.07 ;
      RECT 110.57 365.59 116.41 365.75 ;
      RECT 110.57 362.36 113.2 365.22 ;
      RECT 105.98 364.23 109.06 365.19 ;
      RECT 110.57 364.97 116.41 365.13 ;
      RECT 110.57 364.65 116.41 364.81 ;
      RECT 115.35 364.03 115.51 364.81 ;
      RECT 105.98 362.13 109.21 363.09 ;
      RECT 105.98 362.36 115.11 362.92 ;
      RECT 105.97 362.53 116.41 362.69 ;
      RECT 115.84 361.88 116.41 362.04 ;
      RECT 105.98 360.83 109.21 361.79 ;
      RECT 105.98 361 115.11 361.56 ;
      RECT 105.97 361.23 116.41 361.39 ;
      RECT 110.57 358.7 113.2 361.56 ;
      RECT 115.35 359.11 115.51 359.89 ;
      RECT 105.98 358.73 109.06 359.69 ;
      RECT 110.57 359.11 116.41 359.27 ;
      RECT 110.57 358.79 116.41 358.95 ;
      RECT 110.57 355.56 113.2 358.42 ;
      RECT 110.57 358.17 116.41 358.33 ;
      RECT 102.82 357.42 103.1 358.16 ;
      RECT 106.83 357.56 108.71 358.12 ;
      RECT 105.37 357.56 108.71 358.11 ;
      RECT 103.49 357.46 105.37 358.02 ;
      RECT 110.57 357.85 116.41 358.01 ;
      RECT 115.35 357.23 115.51 358.01 ;
      RECT 102.82 357.47 105.37 358.02 ;
      RECT 109.21 355.56 115.11 356.12 ;
      RECT 109.21 355.73 116.41 355.89 ;
      RECT 115.84 355.08 116.41 355.24 ;
      RECT 106.83 343.96 107.39 355.16 ;
      RECT 105.98 354.03 109.21 354.99 ;
      RECT 105.98 354.2 115.11 354.76 ;
      RECT 105.97 354.43 116.41 354.59 ;
      RECT 110.57 351.9 113.2 354.76 ;
      RECT 115.35 352.31 115.51 353.09 ;
      RECT 105.98 351.93 109.06 352.89 ;
      RECT 110.57 352.31 116.41 352.47 ;
      RECT 110.57 351.99 116.41 352.15 ;
      RECT 110.57 348.76 113.2 351.62 ;
      RECT 105.98 350.63 109.06 351.59 ;
      RECT 110.57 351.37 116.41 351.53 ;
      RECT 110.57 351.05 116.41 351.21 ;
      RECT 115.35 350.43 115.51 351.21 ;
      RECT 105.98 348.53 109.21 349.49 ;
      RECT 105.98 348.76 115.11 349.32 ;
      RECT 105.97 348.93 116.41 349.09 ;
      RECT 115.84 348.28 116.41 348.44 ;
      RECT 105.98 347.23 109.21 348.19 ;
      RECT 105.98 347.4 115.11 347.96 ;
      RECT 105.97 347.63 116.41 347.79 ;
      RECT 110.57 345.1 113.2 347.96 ;
      RECT 115.35 345.51 115.51 346.29 ;
      RECT 105.98 345.13 109.06 346.09 ;
      RECT 110.57 345.51 116.41 345.67 ;
      RECT 110.57 345.19 116.41 345.35 ;
      RECT 110.57 341.96 113.2 344.82 ;
      RECT 110.57 344.57 116.41 344.73 ;
      RECT 102.82 343.82 103.1 344.56 ;
      RECT 106.83 343.96 108.71 344.52 ;
      RECT 105.37 343.96 108.71 344.51 ;
      RECT 103.49 343.86 105.37 344.42 ;
      RECT 110.57 344.25 116.41 344.41 ;
      RECT 115.35 343.63 115.51 344.41 ;
      RECT 102.82 343.87 105.37 344.42 ;
      RECT 109.21 341.96 115.11 342.52 ;
      RECT 109.21 342.13 116.41 342.29 ;
      RECT 115.84 341.48 116.41 341.64 ;
      RECT 106.83 330.36 107.39 341.56 ;
      RECT 105.98 340.43 109.21 341.39 ;
      RECT 105.98 340.6 115.11 341.16 ;
      RECT 105.97 340.83 116.41 340.99 ;
      RECT 110.57 338.3 113.2 341.16 ;
      RECT 115.35 338.71 115.51 339.49 ;
      RECT 105.98 338.33 109.06 339.29 ;
      RECT 110.57 338.71 116.41 338.87 ;
      RECT 110.57 338.39 116.41 338.55 ;
      RECT 110.57 335.16 113.2 338.02 ;
      RECT 105.98 337.03 109.06 337.99 ;
      RECT 110.57 337.77 116.41 337.93 ;
      RECT 110.57 337.45 116.41 337.61 ;
      RECT 115.35 336.83 115.51 337.61 ;
      RECT 105.98 334.93 109.21 335.89 ;
      RECT 105.98 335.16 115.11 335.72 ;
      RECT 105.97 335.33 116.41 335.49 ;
      RECT 115.84 334.68 116.41 334.84 ;
      RECT 105.98 333.63 109.21 334.59 ;
      RECT 105.98 333.8 115.11 334.36 ;
      RECT 105.97 334.03 116.41 334.19 ;
      RECT 110.57 331.5 113.2 334.36 ;
      RECT 115.35 331.91 115.51 332.69 ;
      RECT 105.98 331.53 109.06 332.49 ;
      RECT 110.57 331.91 116.41 332.07 ;
      RECT 110.57 331.59 116.41 331.75 ;
      RECT 110.57 328.36 113.2 331.22 ;
      RECT 110.57 330.97 116.41 331.13 ;
      RECT 102.82 330.22 103.1 330.96 ;
      RECT 106.83 330.36 108.71 330.92 ;
      RECT 105.37 330.36 108.71 330.91 ;
      RECT 103.49 330.26 105.37 330.82 ;
      RECT 110.57 330.65 116.41 330.81 ;
      RECT 115.35 330.03 115.51 330.81 ;
      RECT 102.82 330.27 105.37 330.82 ;
      RECT 109.21 328.36 115.11 328.92 ;
      RECT 109.21 328.53 116.41 328.69 ;
      RECT 115.84 327.88 116.41 328.04 ;
      RECT 106.83 316.76 107.39 327.96 ;
      RECT 105.98 326.83 109.21 327.79 ;
      RECT 105.98 327 115.11 327.56 ;
      RECT 105.97 327.23 116.41 327.39 ;
      RECT 110.57 324.7 113.2 327.56 ;
      RECT 115.35 325.11 115.51 325.89 ;
      RECT 105.98 324.73 109.06 325.69 ;
      RECT 110.57 325.11 116.41 325.27 ;
      RECT 110.57 324.79 116.41 324.95 ;
      RECT 110.57 321.56 113.2 324.42 ;
      RECT 105.98 323.43 109.06 324.39 ;
      RECT 110.57 324.17 116.41 324.33 ;
      RECT 110.57 323.85 116.41 324.01 ;
      RECT 115.35 323.23 115.51 324.01 ;
      RECT 105.98 321.33 109.21 322.29 ;
      RECT 105.98 321.56 115.11 322.12 ;
      RECT 105.97 321.73 116.41 321.89 ;
      RECT 115.84 321.08 116.41 321.24 ;
      RECT 105.98 320.03 109.21 320.99 ;
      RECT 105.98 320.2 115.11 320.76 ;
      RECT 105.97 320.43 116.41 320.59 ;
      RECT 110.57 317.9 113.2 320.76 ;
      RECT 115.35 318.31 115.51 319.09 ;
      RECT 105.98 317.93 109.06 318.89 ;
      RECT 110.57 318.31 116.41 318.47 ;
      RECT 110.57 317.99 116.41 318.15 ;
      RECT 110.57 314.76 113.2 317.62 ;
      RECT 110.57 317.37 116.41 317.53 ;
      RECT 102.82 316.62 103.1 317.36 ;
      RECT 106.83 316.76 108.71 317.32 ;
      RECT 105.37 316.76 108.71 317.31 ;
      RECT 103.49 316.66 105.37 317.22 ;
      RECT 110.57 317.05 116.41 317.21 ;
      RECT 115.35 316.43 115.51 317.21 ;
      RECT 102.82 316.67 105.37 317.22 ;
      RECT 109.21 314.76 115.11 315.32 ;
      RECT 109.21 314.93 116.41 315.09 ;
      RECT 115.84 314.28 116.41 314.44 ;
      RECT 106.83 303.16 107.39 314.36 ;
      RECT 105.98 313.23 109.21 314.19 ;
      RECT 105.98 313.4 115.11 313.96 ;
      RECT 105.97 313.63 116.41 313.79 ;
      RECT 110.57 311.1 113.2 313.96 ;
      RECT 115.35 311.51 115.51 312.29 ;
      RECT 105.98 311.13 109.06 312.09 ;
      RECT 110.57 311.51 116.41 311.67 ;
      RECT 110.57 311.19 116.41 311.35 ;
      RECT 110.57 307.96 113.2 310.82 ;
      RECT 105.98 309.83 109.06 310.79 ;
      RECT 110.57 310.57 116.41 310.73 ;
      RECT 110.57 310.25 116.41 310.41 ;
      RECT 115.35 309.63 115.51 310.41 ;
      RECT 105.98 307.73 109.21 308.69 ;
      RECT 105.98 307.96 115.11 308.52 ;
      RECT 105.97 308.13 116.41 308.29 ;
      RECT 115.84 307.48 116.41 307.64 ;
      RECT 105.98 306.43 109.21 307.39 ;
      RECT 105.98 306.6 115.11 307.16 ;
      RECT 105.97 306.83 116.41 306.99 ;
      RECT 110.57 304.3 113.2 307.16 ;
      RECT 115.35 304.71 115.51 305.49 ;
      RECT 105.98 304.33 109.06 305.29 ;
      RECT 110.57 304.71 116.41 304.87 ;
      RECT 110.57 304.39 116.41 304.55 ;
      RECT 110.57 301.16 113.2 304.02 ;
      RECT 110.57 303.77 116.41 303.93 ;
      RECT 102.82 303.02 103.1 303.76 ;
      RECT 106.83 303.16 108.71 303.72 ;
      RECT 105.37 303.16 108.71 303.71 ;
      RECT 103.49 303.06 105.37 303.62 ;
      RECT 110.57 303.45 116.41 303.61 ;
      RECT 115.35 302.83 115.51 303.61 ;
      RECT 102.82 303.07 105.37 303.62 ;
      RECT 109.21 301.16 115.11 301.72 ;
      RECT 109.21 301.33 116.41 301.49 ;
      RECT 115.84 300.68 116.41 300.84 ;
      RECT 106.83 289.56 107.39 300.76 ;
      RECT 105.98 299.63 109.21 300.59 ;
      RECT 105.98 299.8 115.11 300.36 ;
      RECT 105.97 300.03 116.41 300.19 ;
      RECT 110.57 297.5 113.2 300.36 ;
      RECT 115.35 297.91 115.51 298.69 ;
      RECT 105.98 297.53 109.06 298.49 ;
      RECT 110.57 297.91 116.41 298.07 ;
      RECT 110.57 297.59 116.41 297.75 ;
      RECT 110.57 294.36 113.2 297.22 ;
      RECT 105.98 296.23 109.06 297.19 ;
      RECT 110.57 296.97 116.41 297.13 ;
      RECT 110.57 296.65 116.41 296.81 ;
      RECT 115.35 296.03 115.51 296.81 ;
      RECT 105.98 294.13 109.21 295.09 ;
      RECT 105.98 294.36 115.11 294.92 ;
      RECT 105.97 294.53 116.41 294.69 ;
      RECT 115.84 293.88 116.41 294.04 ;
      RECT 105.98 292.83 109.21 293.79 ;
      RECT 105.98 293 115.11 293.56 ;
      RECT 105.97 293.23 116.41 293.39 ;
      RECT 110.57 290.7 113.2 293.56 ;
      RECT 115.35 291.11 115.51 291.89 ;
      RECT 105.98 290.73 109.06 291.69 ;
      RECT 110.57 291.11 116.41 291.27 ;
      RECT 110.57 290.79 116.41 290.95 ;
      RECT 110.57 287.56 113.2 290.42 ;
      RECT 110.57 290.17 116.41 290.33 ;
      RECT 102.82 289.42 103.1 290.16 ;
      RECT 105.37 289.56 108.71 290.12 ;
      RECT 103.49 289.46 105.37 290.02 ;
      RECT 110.57 289.85 116.41 290.01 ;
      RECT 115.35 289.23 115.51 290.01 ;
      RECT 102.82 289.47 105.37 290.02 ;
      RECT 109.21 287.56 115.11 288.12 ;
      RECT 109.21 287.73 116.41 287.89 ;
      RECT 115.84 287.08 116.41 287.24 ;
      RECT 106.83 275.96 107.39 287.16 ;
      RECT 105.98 286.03 109.21 286.99 ;
      RECT 105.98 286.2 115.11 286.76 ;
      RECT 105.97 286.43 116.41 286.59 ;
      RECT 110.57 283.9 113.2 286.76 ;
      RECT 115.35 284.31 115.51 285.09 ;
      RECT 105.98 283.93 109.06 284.89 ;
      RECT 110.57 284.31 116.41 284.47 ;
      RECT 110.57 283.99 116.41 284.15 ;
      RECT 110.57 280.76 113.2 283.62 ;
      RECT 105.98 282.63 109.06 283.59 ;
      RECT 110.57 283.37 116.41 283.53 ;
      RECT 110.57 283.05 116.41 283.21 ;
      RECT 115.35 282.43 115.51 283.21 ;
      RECT 105.98 280.53 109.21 281.49 ;
      RECT 105.98 280.76 115.11 281.32 ;
      RECT 105.97 280.93 116.41 281.09 ;
      RECT 115.84 280.28 116.41 280.44 ;
      RECT 105.98 279.23 109.21 280.19 ;
      RECT 105.98 279.4 115.11 279.96 ;
      RECT 105.97 279.63 116.41 279.79 ;
      RECT 110.57 277.1 113.2 279.96 ;
      RECT 115.35 277.51 115.51 278.29 ;
      RECT 105.98 277.13 109.06 278.09 ;
      RECT 110.57 277.51 116.41 277.67 ;
      RECT 110.57 277.19 116.41 277.35 ;
      RECT 110.57 273.96 113.2 276.82 ;
      RECT 110.57 276.57 116.41 276.73 ;
      RECT 102.82 275.82 103.1 276.56 ;
      RECT 106.83 275.96 108.71 276.52 ;
      RECT 105.37 275.96 108.71 276.51 ;
      RECT 103.49 275.86 105.37 276.42 ;
      RECT 110.57 276.25 116.41 276.41 ;
      RECT 115.35 275.63 115.51 276.41 ;
      RECT 102.82 275.87 105.37 276.42 ;
      RECT 109.21 273.96 115.11 274.52 ;
      RECT 109.21 274.13 116.41 274.29 ;
      RECT 115.84 273.48 116.41 273.64 ;
      RECT 106.83 262.36 107.39 273.56 ;
      RECT 105.98 272.43 109.21 273.39 ;
      RECT 105.98 272.6 115.11 273.16 ;
      RECT 105.97 272.83 116.41 272.99 ;
      RECT 110.57 270.3 113.2 273.16 ;
      RECT 115.35 270.71 115.51 271.49 ;
      RECT 105.98 270.33 109.06 271.29 ;
      RECT 110.57 270.71 116.41 270.87 ;
      RECT 110.57 270.39 116.41 270.55 ;
      RECT 110.57 267.16 113.2 270.02 ;
      RECT 105.98 269.03 109.06 269.99 ;
      RECT 110.57 269.77 116.41 269.93 ;
      RECT 110.57 269.45 116.41 269.61 ;
      RECT 115.35 268.83 115.51 269.61 ;
      RECT 105.98 266.93 109.21 267.89 ;
      RECT 105.98 267.16 115.11 267.72 ;
      RECT 105.97 267.33 116.41 267.49 ;
      RECT 115.84 266.68 116.41 266.84 ;
      RECT 105.98 265.63 109.21 266.59 ;
      RECT 105.98 265.8 115.11 266.36 ;
      RECT 105.97 266.03 116.41 266.19 ;
      RECT 110.57 263.5 113.2 266.36 ;
      RECT 115.35 263.91 115.51 264.69 ;
      RECT 105.98 263.53 109.06 264.49 ;
      RECT 110.57 263.91 116.41 264.07 ;
      RECT 110.57 263.59 116.41 263.75 ;
      RECT 110.57 260.36 113.2 263.22 ;
      RECT 110.57 262.97 116.41 263.13 ;
      RECT 102.82 262.22 103.1 262.96 ;
      RECT 106.83 262.36 108.71 262.92 ;
      RECT 105.37 262.36 108.71 262.91 ;
      RECT 103.49 262.26 105.37 262.82 ;
      RECT 110.57 262.65 116.41 262.81 ;
      RECT 115.35 262.03 115.51 262.81 ;
      RECT 102.82 262.27 105.37 262.82 ;
      RECT 109.21 260.36 115.11 260.92 ;
      RECT 109.21 260.53 116.41 260.69 ;
      RECT 115.84 259.88 116.41 260.04 ;
      RECT 106.83 248.76 107.39 259.96 ;
      RECT 105.98 258.83 109.21 259.79 ;
      RECT 105.98 259 115.11 259.56 ;
      RECT 105.97 259.23 116.41 259.39 ;
      RECT 110.57 256.7 113.2 259.56 ;
      RECT 115.35 257.11 115.51 257.89 ;
      RECT 105.98 256.73 109.06 257.69 ;
      RECT 110.57 257.11 116.41 257.27 ;
      RECT 110.57 256.79 116.41 256.95 ;
      RECT 110.57 253.56 113.2 256.42 ;
      RECT 105.98 255.43 109.06 256.39 ;
      RECT 110.57 256.17 116.41 256.33 ;
      RECT 110.57 255.85 116.41 256.01 ;
      RECT 115.35 255.23 115.51 256.01 ;
      RECT 105.98 253.33 109.21 254.29 ;
      RECT 105.98 253.56 115.11 254.12 ;
      RECT 105.97 253.73 116.41 253.89 ;
      RECT 115.84 253.08 116.41 253.24 ;
      RECT 105.98 252.03 109.21 252.99 ;
      RECT 105.98 252.2 115.11 252.76 ;
      RECT 105.97 252.43 116.41 252.59 ;
      RECT 110.57 249.9 113.2 252.76 ;
      RECT 115.35 250.31 115.51 251.09 ;
      RECT 105.98 249.93 109.06 250.89 ;
      RECT 110.57 250.31 116.41 250.47 ;
      RECT 110.57 249.99 116.41 250.15 ;
      RECT 110.57 246.76 113.2 249.62 ;
      RECT 110.57 249.37 116.41 249.53 ;
      RECT 102.82 248.62 103.1 249.36 ;
      RECT 106.83 248.76 108.71 249.32 ;
      RECT 105.37 248.76 108.71 249.31 ;
      RECT 103.49 248.66 105.37 249.22 ;
      RECT 110.57 249.05 116.41 249.21 ;
      RECT 115.35 248.43 115.51 249.21 ;
      RECT 102.82 248.67 105.37 249.22 ;
      RECT 109.21 246.76 115.11 247.32 ;
      RECT 109.21 246.93 116.41 247.09 ;
      RECT 115.84 246.28 116.41 246.44 ;
      RECT 106.83 235.16 107.39 246.36 ;
      RECT 105.98 245.23 109.21 246.19 ;
      RECT 105.98 245.4 115.11 245.96 ;
      RECT 105.97 245.63 116.41 245.79 ;
      RECT 110.57 243.1 113.2 245.96 ;
      RECT 115.35 243.51 115.51 244.29 ;
      RECT 105.98 243.13 109.06 244.09 ;
      RECT 110.57 243.51 116.41 243.67 ;
      RECT 110.57 243.19 116.41 243.35 ;
      RECT 110.57 239.96 113.2 242.82 ;
      RECT 105.98 241.83 109.06 242.79 ;
      RECT 110.57 242.57 116.41 242.73 ;
      RECT 110.57 242.25 116.41 242.41 ;
      RECT 115.35 241.63 115.51 242.41 ;
      RECT 105.98 239.73 109.21 240.69 ;
      RECT 105.98 239.96 115.11 240.52 ;
      RECT 105.97 240.13 116.41 240.29 ;
      RECT 115.84 239.48 116.41 239.64 ;
      RECT 105.98 238.43 109.21 239.39 ;
      RECT 105.98 238.6 115.11 239.16 ;
      RECT 105.97 238.83 116.41 238.99 ;
      RECT 110.57 236.3 113.2 239.16 ;
      RECT 115.35 236.71 115.51 237.49 ;
      RECT 105.98 236.33 109.06 237.29 ;
      RECT 110.57 236.71 116.41 236.87 ;
      RECT 110.57 236.39 116.41 236.55 ;
      RECT 110.57 233.16 113.2 236.02 ;
      RECT 110.57 235.77 116.41 235.93 ;
      RECT 102.82 235.02 103.1 235.76 ;
      RECT 106.83 235.16 108.71 235.72 ;
      RECT 105.37 235.16 108.71 235.71 ;
      RECT 103.49 235.06 105.37 235.62 ;
      RECT 110.57 235.45 116.41 235.61 ;
      RECT 115.35 234.83 115.51 235.61 ;
      RECT 102.82 235.07 105.37 235.62 ;
      RECT 109.21 233.16 115.11 233.72 ;
      RECT 109.21 233.33 116.41 233.49 ;
      RECT 115.84 232.68 116.41 232.84 ;
      RECT 106.83 221.56 107.39 232.76 ;
      RECT 105.98 231.63 109.21 232.59 ;
      RECT 105.98 231.8 115.11 232.36 ;
      RECT 105.97 232.03 116.41 232.19 ;
      RECT 110.57 229.5 113.2 232.36 ;
      RECT 115.35 229.91 115.51 230.69 ;
      RECT 105.98 229.53 109.06 230.49 ;
      RECT 110.57 229.91 116.41 230.07 ;
      RECT 110.57 229.59 116.41 229.75 ;
      RECT 110.57 226.36 113.2 229.22 ;
      RECT 105.98 228.23 109.06 229.19 ;
      RECT 110.57 228.97 116.41 229.13 ;
      RECT 110.57 228.65 116.41 228.81 ;
      RECT 115.35 228.03 115.51 228.81 ;
      RECT 105.98 226.13 109.21 227.09 ;
      RECT 105.98 226.36 115.11 226.92 ;
      RECT 105.97 226.53 116.41 226.69 ;
      RECT 115.84 225.88 116.41 226.04 ;
      RECT 105.98 224.83 109.21 225.79 ;
      RECT 105.98 225 115.11 225.56 ;
      RECT 105.97 225.23 116.41 225.39 ;
      RECT 110.57 222.7 113.2 225.56 ;
      RECT 115.35 223.11 115.51 223.89 ;
      RECT 105.98 222.73 109.06 223.69 ;
      RECT 110.57 223.11 116.41 223.27 ;
      RECT 110.57 222.79 116.41 222.95 ;
      RECT 110.57 219.56 113.2 222.42 ;
      RECT 110.57 222.17 116.41 222.33 ;
      RECT 102.82 221.42 103.1 222.16 ;
      RECT 106.83 221.56 108.71 222.12 ;
      RECT 105.37 221.56 108.71 222.11 ;
      RECT 103.49 221.46 105.37 222.02 ;
      RECT 110.57 221.85 116.41 222.01 ;
      RECT 115.35 221.23 115.51 222.01 ;
      RECT 102.82 221.47 105.37 222.02 ;
      RECT 109.21 219.56 115.11 220.12 ;
      RECT 109.21 219.73 116.41 219.89 ;
      RECT 115.84 219.08 116.41 219.24 ;
      RECT 115.84 212.28 116.41 212.44 ;
      RECT 110.57 205.96 113.2 208.82 ;
      RECT 110.57 208.57 116.41 208.73 ;
      RECT 110.57 208.25 116.41 208.41 ;
      RECT 115.35 207.63 115.51 208.41 ;
      RECT 109.21 205.96 115.11 206.52 ;
      RECT 109.21 206.13 116.41 206.29 ;
      RECT 110.57 192.36 113.2 195.22 ;
      RECT 110.57 194.97 116.41 195.13 ;
      RECT 110.57 194.65 116.41 194.81 ;
      RECT 115.35 194.03 115.51 194.81 ;
      RECT 109.21 192.36 115.11 192.92 ;
      RECT 109.21 192.53 116.41 192.69 ;
      RECT 110.57 178.76 113.2 181.62 ;
      RECT 110.57 181.37 116.41 181.53 ;
      RECT 110.57 181.05 116.41 181.21 ;
      RECT 115.35 180.43 115.51 181.21 ;
      RECT 109.21 178.76 115.11 179.32 ;
      RECT 109.21 178.93 116.41 179.09 ;
      RECT 110.57 165.16 113.2 168.02 ;
      RECT 110.57 167.77 116.41 167.93 ;
      RECT 110.57 167.45 116.41 167.61 ;
      RECT 115.35 166.83 115.51 167.61 ;
      RECT 109.21 165.16 115.11 165.72 ;
      RECT 109.21 165.33 116.41 165.49 ;
      RECT 110.57 151.56 113.2 154.42 ;
      RECT 110.57 154.17 116.41 154.33 ;
      RECT 110.57 153.85 116.41 154.01 ;
      RECT 115.35 153.23 115.51 154.01 ;
      RECT 109.21 151.56 115.11 152.12 ;
      RECT 109.21 151.73 116.41 151.89 ;
      RECT 110.57 137.96 113.2 140.82 ;
      RECT 110.57 140.57 116.41 140.73 ;
      RECT 110.57 140.25 116.41 140.41 ;
      RECT 115.35 139.63 115.51 140.41 ;
      RECT 109.21 137.96 115.11 138.52 ;
      RECT 109.21 138.13 116.41 138.29 ;
      RECT 115.84 69.48 116.41 69.64 ;
      RECT 115.93 31.49 116.09 32.02 ;
      RECT 115.47 31.49 116.55 31.65 ;
      RECT 116.39 27.38 116.55 31.65 ;
      RECT 115.47 27.38 115.63 31.65 ;
      RECT 115.47 27.38 116.55 27.54 ;
      RECT 115.93 26.91 116.09 27.54 ;
      RECT 115.47 51.06 116.55 55.29 ;
      RECT 115.93 50.27 116.09 55.29 ;
      RECT 116.29 49.92 116.45 50.9 ;
      RECT 115.57 49.92 115.73 50.9 ;
      RECT 115.57 49.92 116.45 50.08 ;
      RECT 115.93 45.65 116.09 50.08 ;
      RECT 110.57 69.96 113.2 72.82 ;
      RECT 110.57 72.57 116.25 72.73 ;
      RECT 110.57 72.25 116.25 72.41 ;
      RECT 115.35 71.63 115.51 72.41 ;
      RECT 109.21 69.96 115.11 70.52 ;
      RECT 109.21 70.13 116.25 70.29 ;
      RECT 106.83 72.96 107.39 83.16 ;
      RECT 105.98 82.03 109.21 82.99 ;
      RECT 105.98 82.2 115.11 82.76 ;
      RECT 105.97 82.43 116.25 82.59 ;
      RECT 110.57 79.9 113.2 82.76 ;
      RECT 115.35 80.31 115.51 81.09 ;
      RECT 105.98 79.93 109.06 80.89 ;
      RECT 110.57 80.31 116.25 80.47 ;
      RECT 110.57 79.99 116.25 80.15 ;
      RECT 110.57 76.76 113.2 79.62 ;
      RECT 105.98 78.63 109.06 79.59 ;
      RECT 110.57 79.37 116.25 79.53 ;
      RECT 110.57 79.05 116.25 79.21 ;
      RECT 115.35 78.43 115.51 79.21 ;
      RECT 105.98 76.53 109.21 77.49 ;
      RECT 105.98 76.76 115.11 77.32 ;
      RECT 105.97 76.93 116.25 77.09 ;
      RECT 105.98 75.23 109.21 76.19 ;
      RECT 105.98 75.4 115.11 75.96 ;
      RECT 105.97 75.63 116.25 75.79 ;
      RECT 110.57 73.1 113.2 75.96 ;
      RECT 115.35 73.51 115.51 74.29 ;
      RECT 105.98 73.13 109.06 74.09 ;
      RECT 110.57 73.51 116.25 73.67 ;
      RECT 110.57 73.19 116.25 73.35 ;
      RECT 110.57 83.56 113.2 86.42 ;
      RECT 110.57 86.17 116.25 86.33 ;
      RECT 110.57 85.85 116.25 86.01 ;
      RECT 115.35 85.23 115.51 86.01 ;
      RECT 109.21 83.56 115.11 84.12 ;
      RECT 109.21 83.73 116.25 83.89 ;
      RECT 106.83 85.56 107.39 96.76 ;
      RECT 105.98 95.63 109.21 96.59 ;
      RECT 105.98 95.8 115.11 96.36 ;
      RECT 105.97 96.03 116.25 96.19 ;
      RECT 110.57 93.5 113.2 96.36 ;
      RECT 115.35 93.91 115.51 94.69 ;
      RECT 105.98 93.53 109.06 94.49 ;
      RECT 110.57 93.91 116.25 94.07 ;
      RECT 110.57 93.59 116.25 93.75 ;
      RECT 110.57 90.36 113.2 93.22 ;
      RECT 105.98 92.23 109.06 93.19 ;
      RECT 110.57 92.97 116.25 93.13 ;
      RECT 110.57 92.65 116.25 92.81 ;
      RECT 115.35 92.03 115.51 92.81 ;
      RECT 105.98 90.13 109.21 91.09 ;
      RECT 105.98 90.36 115.11 90.92 ;
      RECT 105.97 90.53 116.25 90.69 ;
      RECT 105.98 88.83 109.21 89.79 ;
      RECT 105.98 89 115.11 89.56 ;
      RECT 105.97 89.23 116.25 89.39 ;
      RECT 110.57 86.7 113.2 89.56 ;
      RECT 115.35 87.11 115.51 87.89 ;
      RECT 105.98 86.73 109.06 87.69 ;
      RECT 110.57 87.11 116.25 87.27 ;
      RECT 110.57 86.79 116.25 86.95 ;
      RECT 102.82 85.42 103.1 86.16 ;
      RECT 106.83 85.56 108.71 86.12 ;
      RECT 105.37 85.56 108.71 86.11 ;
      RECT 103.49 85.46 105.37 86.02 ;
      RECT 102.82 85.47 105.37 86.02 ;
      RECT 110.57 97.16 113.2 100.02 ;
      RECT 110.57 99.77 116.25 99.93 ;
      RECT 110.57 99.45 116.25 99.61 ;
      RECT 115.35 98.83 115.51 99.61 ;
      RECT 109.21 97.16 115.11 97.72 ;
      RECT 109.21 97.33 116.25 97.49 ;
      RECT 106.83 99.16 107.39 110.36 ;
      RECT 105.98 109.23 109.21 110.19 ;
      RECT 105.98 109.4 115.11 109.96 ;
      RECT 105.97 109.63 116.25 109.79 ;
      RECT 110.57 107.1 113.2 109.96 ;
      RECT 115.35 107.51 115.51 108.29 ;
      RECT 105.98 107.13 109.06 108.09 ;
      RECT 110.57 107.51 116.25 107.67 ;
      RECT 110.57 107.19 116.25 107.35 ;
      RECT 110.57 103.96 113.2 106.82 ;
      RECT 105.98 105.83 109.06 106.79 ;
      RECT 110.57 106.57 116.25 106.73 ;
      RECT 110.57 106.25 116.25 106.41 ;
      RECT 115.35 105.63 115.51 106.41 ;
      RECT 105.98 103.73 109.21 104.69 ;
      RECT 105.98 103.96 115.11 104.52 ;
      RECT 105.97 104.13 116.25 104.29 ;
      RECT 105.98 102.43 109.21 103.39 ;
      RECT 105.98 102.6 115.11 103.16 ;
      RECT 105.97 102.83 116.25 102.99 ;
      RECT 110.57 100.3 113.2 103.16 ;
      RECT 115.35 100.71 115.51 101.49 ;
      RECT 105.98 100.33 109.06 101.29 ;
      RECT 110.57 100.71 116.25 100.87 ;
      RECT 110.57 100.39 116.25 100.55 ;
      RECT 102.82 99.02 103.1 99.76 ;
      RECT 106.83 99.16 108.71 99.72 ;
      RECT 105.37 99.16 108.71 99.71 ;
      RECT 103.49 99.06 105.37 99.62 ;
      RECT 102.82 99.07 105.37 99.62 ;
      RECT 110.57 110.76 113.2 113.62 ;
      RECT 110.57 113.37 116.25 113.53 ;
      RECT 110.57 113.05 116.25 113.21 ;
      RECT 115.35 112.43 115.51 113.21 ;
      RECT 109.21 110.76 115.11 111.32 ;
      RECT 109.21 110.93 116.25 111.09 ;
      RECT 106.83 112.76 107.39 123.96 ;
      RECT 105.98 122.83 109.21 123.79 ;
      RECT 105.98 123 115.11 123.56 ;
      RECT 105.97 123.23 116.25 123.39 ;
      RECT 110.57 120.7 113.2 123.56 ;
      RECT 115.35 121.11 115.51 121.89 ;
      RECT 105.98 120.73 109.06 121.69 ;
      RECT 110.57 121.11 116.25 121.27 ;
      RECT 110.57 120.79 116.25 120.95 ;
      RECT 110.57 117.56 113.2 120.42 ;
      RECT 105.98 119.43 109.06 120.39 ;
      RECT 110.57 120.17 116.25 120.33 ;
      RECT 110.57 119.85 116.25 120.01 ;
      RECT 115.35 119.23 115.51 120.01 ;
      RECT 105.98 117.33 109.21 118.29 ;
      RECT 105.98 117.56 115.11 118.12 ;
      RECT 105.97 117.73 116.25 117.89 ;
      RECT 105.98 116.03 109.21 116.99 ;
      RECT 105.98 116.2 115.11 116.76 ;
      RECT 105.97 116.43 116.25 116.59 ;
      RECT 110.57 113.9 113.2 116.76 ;
      RECT 115.35 114.31 115.51 115.09 ;
      RECT 105.98 113.93 109.06 114.89 ;
      RECT 110.57 114.31 116.25 114.47 ;
      RECT 110.57 113.99 116.25 114.15 ;
      RECT 102.82 112.62 103.1 113.36 ;
      RECT 106.83 112.76 108.71 113.32 ;
      RECT 105.37 112.76 108.71 113.31 ;
      RECT 103.49 112.66 105.37 113.22 ;
      RECT 102.82 112.67 105.37 113.22 ;
      RECT 110.57 124.36 113.2 127.22 ;
      RECT 110.57 126.97 116.25 127.13 ;
      RECT 110.57 126.65 116.25 126.81 ;
      RECT 115.35 126.03 115.51 126.81 ;
      RECT 109.21 124.36 115.11 124.92 ;
      RECT 109.21 124.53 116.25 124.69 ;
      RECT 106.83 126.36 107.39 137.56 ;
      RECT 105.98 136.43 109.21 137.39 ;
      RECT 105.98 136.6 115.11 137.16 ;
      RECT 105.97 136.83 116.25 136.99 ;
      RECT 110.57 134.3 113.2 137.16 ;
      RECT 115.35 134.71 115.51 135.49 ;
      RECT 105.98 134.33 109.06 135.29 ;
      RECT 110.57 134.71 116.25 134.87 ;
      RECT 110.57 134.39 116.25 134.55 ;
      RECT 110.57 131.16 113.2 134.02 ;
      RECT 105.98 133.03 109.06 133.99 ;
      RECT 110.57 133.77 116.25 133.93 ;
      RECT 110.57 133.45 116.25 133.61 ;
      RECT 115.35 132.83 115.51 133.61 ;
      RECT 105.98 130.93 109.21 131.89 ;
      RECT 105.98 131.16 115.11 131.72 ;
      RECT 105.97 131.33 116.25 131.49 ;
      RECT 105.98 129.63 109.21 130.59 ;
      RECT 105.98 129.8 115.11 130.36 ;
      RECT 105.97 130.03 116.25 130.19 ;
      RECT 110.57 127.5 113.2 130.36 ;
      RECT 115.35 127.91 115.51 128.69 ;
      RECT 105.98 127.53 109.06 128.49 ;
      RECT 110.57 127.91 116.25 128.07 ;
      RECT 110.57 127.59 116.25 127.75 ;
      RECT 102.82 126.22 103.1 126.96 ;
      RECT 106.83 126.36 108.71 126.92 ;
      RECT 105.37 126.36 108.71 126.91 ;
      RECT 103.49 126.26 105.37 126.82 ;
      RECT 102.82 126.27 105.37 126.82 ;
      RECT 106.83 139.96 107.39 151.16 ;
      RECT 105.98 150.03 109.21 150.99 ;
      RECT 105.98 150.2 115.11 150.76 ;
      RECT 105.97 150.43 116.25 150.59 ;
      RECT 110.57 147.9 113.2 150.76 ;
      RECT 115.35 148.31 115.51 149.09 ;
      RECT 105.98 147.93 109.06 148.89 ;
      RECT 110.57 148.31 116.25 148.47 ;
      RECT 110.57 147.99 116.25 148.15 ;
      RECT 110.57 144.76 113.2 147.62 ;
      RECT 105.98 146.63 109.06 147.59 ;
      RECT 110.57 147.37 116.25 147.53 ;
      RECT 110.57 147.05 116.25 147.21 ;
      RECT 115.35 146.43 115.51 147.21 ;
      RECT 105.98 144.53 109.21 145.49 ;
      RECT 105.98 144.76 115.11 145.32 ;
      RECT 105.97 144.93 116.25 145.09 ;
      RECT 105.98 143.23 109.21 144.19 ;
      RECT 105.98 143.4 115.11 143.96 ;
      RECT 105.97 143.63 116.25 143.79 ;
      RECT 110.57 141.1 113.2 143.96 ;
      RECT 115.35 141.51 115.51 142.29 ;
      RECT 105.98 141.13 109.06 142.09 ;
      RECT 110.57 141.51 116.25 141.67 ;
      RECT 110.57 141.19 116.25 141.35 ;
      RECT 102.82 139.82 103.1 140.56 ;
      RECT 106.83 139.96 108.71 140.52 ;
      RECT 105.37 139.96 108.71 140.51 ;
      RECT 103.49 139.86 105.37 140.42 ;
      RECT 102.82 139.87 105.37 140.42 ;
      RECT 106.83 153.56 107.39 164.76 ;
      RECT 105.98 163.63 109.21 164.59 ;
      RECT 105.98 163.8 115.11 164.36 ;
      RECT 105.97 164.03 116.25 164.19 ;
      RECT 110.57 161.5 113.2 164.36 ;
      RECT 115.35 161.91 115.51 162.69 ;
      RECT 105.98 161.53 109.06 162.49 ;
      RECT 110.57 161.91 116.25 162.07 ;
      RECT 110.57 161.59 116.25 161.75 ;
      RECT 110.57 158.36 113.2 161.22 ;
      RECT 105.98 160.23 109.06 161.19 ;
      RECT 110.57 160.97 116.25 161.13 ;
      RECT 110.57 160.65 116.25 160.81 ;
      RECT 115.35 160.03 115.51 160.81 ;
      RECT 105.98 158.13 109.21 159.09 ;
      RECT 105.98 158.36 115.11 158.92 ;
      RECT 105.97 158.53 116.25 158.69 ;
      RECT 105.98 156.83 109.21 157.79 ;
      RECT 105.98 157 115.11 157.56 ;
      RECT 105.97 157.23 116.25 157.39 ;
      RECT 110.57 154.7 113.2 157.56 ;
      RECT 115.35 155.11 115.51 155.89 ;
      RECT 105.98 154.73 109.06 155.69 ;
      RECT 110.57 155.11 116.25 155.27 ;
      RECT 110.57 154.79 116.25 154.95 ;
      RECT 102.82 153.42 103.1 154.16 ;
      RECT 106.83 153.56 108.71 154.12 ;
      RECT 105.37 153.56 108.71 154.11 ;
      RECT 103.49 153.46 105.37 154.02 ;
      RECT 102.82 153.47 105.37 154.02 ;
      RECT 106.83 167.16 107.39 178.36 ;
      RECT 105.98 177.23 109.21 178.19 ;
      RECT 105.98 177.4 115.11 177.96 ;
      RECT 105.97 177.63 116.25 177.79 ;
      RECT 110.57 175.1 113.2 177.96 ;
      RECT 115.35 175.51 115.51 176.29 ;
      RECT 105.98 175.13 109.06 176.09 ;
      RECT 110.57 175.51 116.25 175.67 ;
      RECT 110.57 175.19 116.25 175.35 ;
      RECT 110.57 171.96 113.2 174.82 ;
      RECT 105.98 173.83 109.06 174.79 ;
      RECT 110.57 174.57 116.25 174.73 ;
      RECT 110.57 174.25 116.25 174.41 ;
      RECT 115.35 173.63 115.51 174.41 ;
      RECT 105.98 171.73 109.21 172.69 ;
      RECT 105.98 171.96 115.11 172.52 ;
      RECT 105.97 172.13 116.25 172.29 ;
      RECT 105.98 170.43 109.21 171.39 ;
      RECT 105.98 170.6 115.11 171.16 ;
      RECT 105.97 170.83 116.25 170.99 ;
      RECT 110.57 168.3 113.2 171.16 ;
      RECT 115.35 168.71 115.51 169.49 ;
      RECT 105.98 168.33 109.06 169.29 ;
      RECT 110.57 168.71 116.25 168.87 ;
      RECT 110.57 168.39 116.25 168.55 ;
      RECT 102.82 167.02 103.1 167.76 ;
      RECT 106.83 167.16 108.71 167.72 ;
      RECT 105.37 167.16 108.71 167.71 ;
      RECT 103.49 167.06 105.37 167.62 ;
      RECT 102.82 167.07 105.37 167.62 ;
      RECT 106.83 180.76 107.39 191.96 ;
      RECT 105.98 190.83 109.21 191.79 ;
      RECT 105.98 191 115.11 191.56 ;
      RECT 105.97 191.23 116.25 191.39 ;
      RECT 110.57 188.7 113.2 191.56 ;
      RECT 115.35 189.11 115.51 189.89 ;
      RECT 105.98 188.73 109.06 189.69 ;
      RECT 110.57 189.11 116.25 189.27 ;
      RECT 110.57 188.79 116.25 188.95 ;
      RECT 110.57 185.56 113.2 188.42 ;
      RECT 105.98 187.43 109.06 188.39 ;
      RECT 110.57 188.17 116.25 188.33 ;
      RECT 110.57 187.85 116.25 188.01 ;
      RECT 115.35 187.23 115.51 188.01 ;
      RECT 105.98 185.33 109.21 186.29 ;
      RECT 105.98 185.56 115.11 186.12 ;
      RECT 105.97 185.73 116.25 185.89 ;
      RECT 105.98 184.03 109.21 184.99 ;
      RECT 105.98 184.2 115.11 184.76 ;
      RECT 105.97 184.43 116.25 184.59 ;
      RECT 110.57 181.9 113.2 184.76 ;
      RECT 115.35 182.31 115.51 183.09 ;
      RECT 105.98 181.93 109.06 182.89 ;
      RECT 110.57 182.31 116.25 182.47 ;
      RECT 110.57 181.99 116.25 182.15 ;
      RECT 102.82 180.62 103.1 181.36 ;
      RECT 105.37 180.76 108.71 181.32 ;
      RECT 103.49 180.66 105.37 181.22 ;
      RECT 102.82 180.67 105.37 181.22 ;
      RECT 106.83 194.36 107.39 205.56 ;
      RECT 105.98 204.43 109.21 205.39 ;
      RECT 105.98 204.6 115.11 205.16 ;
      RECT 105.97 204.83 116.25 204.99 ;
      RECT 110.57 202.3 113.2 205.16 ;
      RECT 115.35 202.71 115.51 203.49 ;
      RECT 105.98 202.33 109.06 203.29 ;
      RECT 110.57 202.71 116.25 202.87 ;
      RECT 110.57 202.39 116.25 202.55 ;
      RECT 110.57 199.16 113.2 202.02 ;
      RECT 105.98 201.03 109.06 201.99 ;
      RECT 110.57 201.77 116.25 201.93 ;
      RECT 110.57 201.45 116.25 201.61 ;
      RECT 115.35 200.83 115.51 201.61 ;
      RECT 105.98 198.93 109.21 199.89 ;
      RECT 105.98 199.16 115.11 199.72 ;
      RECT 105.97 199.33 116.25 199.49 ;
      RECT 105.98 197.63 109.21 198.59 ;
      RECT 105.98 197.8 115.11 198.36 ;
      RECT 105.97 198.03 116.25 198.19 ;
      RECT 110.57 195.5 113.2 198.36 ;
      RECT 115.35 195.91 115.51 196.69 ;
      RECT 105.98 195.53 109.06 196.49 ;
      RECT 110.57 195.91 116.25 196.07 ;
      RECT 110.57 195.59 116.25 195.75 ;
      RECT 102.82 194.22 103.1 194.96 ;
      RECT 106.83 194.36 108.71 194.92 ;
      RECT 105.37 194.36 108.71 194.91 ;
      RECT 103.49 194.26 105.37 194.82 ;
      RECT 102.82 194.27 105.37 194.82 ;
      RECT 106.83 207.96 107.39 219.16 ;
      RECT 105.98 218.03 109.21 218.99 ;
      RECT 105.98 218.2 115.11 218.76 ;
      RECT 105.97 218.43 116.25 218.59 ;
      RECT 110.57 215.9 113.2 218.76 ;
      RECT 115.35 216.31 115.51 217.09 ;
      RECT 105.98 215.93 109.06 216.89 ;
      RECT 110.57 216.31 116.25 216.47 ;
      RECT 110.57 215.99 116.25 216.15 ;
      RECT 110.57 212.76 113.2 215.62 ;
      RECT 105.98 214.63 109.06 215.59 ;
      RECT 110.57 215.37 116.25 215.53 ;
      RECT 110.57 215.05 116.25 215.21 ;
      RECT 115.35 214.43 115.51 215.21 ;
      RECT 105.98 212.53 109.21 213.49 ;
      RECT 105.98 212.76 115.11 213.32 ;
      RECT 105.97 212.93 116.25 213.09 ;
      RECT 105.98 211.23 109.21 212.19 ;
      RECT 105.98 211.4 115.11 211.96 ;
      RECT 105.97 211.63 116.25 211.79 ;
      RECT 110.57 209.1 113.2 211.96 ;
      RECT 115.35 209.51 115.51 210.29 ;
      RECT 105.98 209.13 109.06 210.09 ;
      RECT 110.57 209.51 116.25 209.67 ;
      RECT 110.57 209.19 116.25 209.35 ;
      RECT 102.82 207.82 103.1 208.56 ;
      RECT 106.83 207.96 108.71 208.52 ;
      RECT 105.37 207.96 108.71 208.51 ;
      RECT 103.49 207.86 105.37 208.42 ;
      RECT 102.82 207.87 105.37 208.42 ;
      RECT 115.85 70.46 116.01 72.05 ;
      RECT 115.13 70.98 116.01 71.14 ;
      RECT 115.85 73.87 116.01 75.46 ;
      RECT 115.13 74.78 116.01 74.94 ;
      RECT 115.85 77.26 116.01 78.85 ;
      RECT 115.13 77.78 116.01 77.94 ;
      RECT 115.85 80.67 116.01 82.26 ;
      RECT 115.13 81.58 116.01 81.74 ;
      RECT 115.85 84.06 116.01 85.65 ;
      RECT 115.13 84.58 116.01 84.74 ;
      RECT 115.85 87.47 116.01 89.06 ;
      RECT 115.13 88.38 116.01 88.54 ;
      RECT 115.85 90.86 116.01 92.45 ;
      RECT 115.13 91.38 116.01 91.54 ;
      RECT 115.85 94.27 116.01 95.86 ;
      RECT 115.13 95.18 116.01 95.34 ;
      RECT 115.85 97.66 116.01 99.25 ;
      RECT 115.13 98.18 116.01 98.34 ;
      RECT 115.85 101.07 116.01 102.66 ;
      RECT 115.13 101.98 116.01 102.14 ;
      RECT 115.85 104.46 116.01 106.05 ;
      RECT 115.13 104.98 116.01 105.14 ;
      RECT 115.85 107.87 116.01 109.46 ;
      RECT 115.13 108.78 116.01 108.94 ;
      RECT 115.85 111.26 116.01 112.85 ;
      RECT 115.13 111.78 116.01 111.94 ;
      RECT 115.85 114.67 116.01 116.26 ;
      RECT 115.13 115.58 116.01 115.74 ;
      RECT 115.85 118.06 116.01 119.65 ;
      RECT 115.13 118.58 116.01 118.74 ;
      RECT 115.85 121.47 116.01 123.06 ;
      RECT 115.13 122.38 116.01 122.54 ;
      RECT 115.85 124.86 116.01 126.45 ;
      RECT 115.13 125.38 116.01 125.54 ;
      RECT 115.85 128.27 116.01 129.86 ;
      RECT 115.13 129.18 116.01 129.34 ;
      RECT 115.85 131.66 116.01 133.25 ;
      RECT 115.13 132.18 116.01 132.34 ;
      RECT 115.85 135.07 116.01 136.66 ;
      RECT 115.13 135.98 116.01 136.14 ;
      RECT 115.85 138.46 116.01 140.05 ;
      RECT 115.13 138.98 116.01 139.14 ;
      RECT 115.85 141.87 116.01 143.46 ;
      RECT 115.13 142.78 116.01 142.94 ;
      RECT 115.85 145.26 116.01 146.85 ;
      RECT 115.13 145.78 116.01 145.94 ;
      RECT 115.85 148.67 116.01 150.26 ;
      RECT 115.13 149.58 116.01 149.74 ;
      RECT 115.85 152.06 116.01 153.65 ;
      RECT 115.13 152.58 116.01 152.74 ;
      RECT 115.85 155.47 116.01 157.06 ;
      RECT 115.13 156.38 116.01 156.54 ;
      RECT 115.85 158.86 116.01 160.45 ;
      RECT 115.13 159.38 116.01 159.54 ;
      RECT 115.85 162.27 116.01 163.86 ;
      RECT 115.13 163.18 116.01 163.34 ;
      RECT 115.85 165.66 116.01 167.25 ;
      RECT 115.13 166.18 116.01 166.34 ;
      RECT 115.85 169.07 116.01 170.66 ;
      RECT 115.13 169.98 116.01 170.14 ;
      RECT 115.85 172.46 116.01 174.05 ;
      RECT 115.13 172.98 116.01 173.14 ;
      RECT 115.85 175.87 116.01 177.46 ;
      RECT 115.13 176.78 116.01 176.94 ;
      RECT 115.85 179.26 116.01 180.85 ;
      RECT 115.13 179.78 116.01 179.94 ;
      RECT 115.85 182.67 116.01 184.26 ;
      RECT 115.13 183.58 116.01 183.74 ;
      RECT 115.85 186.06 116.01 187.65 ;
      RECT 115.13 186.58 116.01 186.74 ;
      RECT 115.85 189.47 116.01 191.06 ;
      RECT 115.13 190.38 116.01 190.54 ;
      RECT 115.85 192.86 116.01 194.45 ;
      RECT 115.13 193.38 116.01 193.54 ;
      RECT 115.85 196.27 116.01 197.86 ;
      RECT 115.13 197.18 116.01 197.34 ;
      RECT 115.85 199.66 116.01 201.25 ;
      RECT 115.13 200.18 116.01 200.34 ;
      RECT 115.85 203.07 116.01 204.66 ;
      RECT 115.13 203.98 116.01 204.14 ;
      RECT 115.85 206.46 116.01 208.05 ;
      RECT 115.13 206.98 116.01 207.14 ;
      RECT 115.85 209.87 116.01 211.46 ;
      RECT 115.13 210.78 116.01 210.94 ;
      RECT 115.85 213.26 116.01 214.85 ;
      RECT 115.13 213.78 116.01 213.94 ;
      RECT 115.85 216.67 116.01 218.26 ;
      RECT 115.13 217.58 116.01 217.74 ;
      RECT 115.85 220.06 116.01 221.65 ;
      RECT 115.13 220.58 116.01 220.74 ;
      RECT 115.85 223.47 116.01 225.06 ;
      RECT 115.13 224.38 116.01 224.54 ;
      RECT 115.85 226.86 116.01 228.45 ;
      RECT 115.13 227.38 116.01 227.54 ;
      RECT 115.85 230.27 116.01 231.86 ;
      RECT 115.13 231.18 116.01 231.34 ;
      RECT 115.85 233.66 116.01 235.25 ;
      RECT 115.13 234.18 116.01 234.34 ;
      RECT 115.85 237.07 116.01 238.66 ;
      RECT 115.13 237.98 116.01 238.14 ;
      RECT 115.85 240.46 116.01 242.05 ;
      RECT 115.13 240.98 116.01 241.14 ;
      RECT 115.85 243.87 116.01 245.46 ;
      RECT 115.13 244.78 116.01 244.94 ;
      RECT 115.85 247.26 116.01 248.85 ;
      RECT 115.13 247.78 116.01 247.94 ;
      RECT 115.85 250.67 116.01 252.26 ;
      RECT 115.13 251.58 116.01 251.74 ;
      RECT 115.85 254.06 116.01 255.65 ;
      RECT 115.13 254.58 116.01 254.74 ;
      RECT 115.85 257.47 116.01 259.06 ;
      RECT 115.13 258.38 116.01 258.54 ;
      RECT 115.85 260.86 116.01 262.45 ;
      RECT 115.13 261.38 116.01 261.54 ;
      RECT 115.85 264.27 116.01 265.86 ;
      RECT 115.13 265.18 116.01 265.34 ;
      RECT 115.85 267.66 116.01 269.25 ;
      RECT 115.13 268.18 116.01 268.34 ;
      RECT 115.85 271.07 116.01 272.66 ;
      RECT 115.13 271.98 116.01 272.14 ;
      RECT 115.85 274.46 116.01 276.05 ;
      RECT 115.13 274.98 116.01 275.14 ;
      RECT 115.85 277.87 116.01 279.46 ;
      RECT 115.13 278.78 116.01 278.94 ;
      RECT 115.85 281.26 116.01 282.85 ;
      RECT 115.13 281.78 116.01 281.94 ;
      RECT 115.85 284.67 116.01 286.26 ;
      RECT 115.13 285.58 116.01 285.74 ;
      RECT 115.85 288.06 116.01 289.65 ;
      RECT 115.13 288.58 116.01 288.74 ;
      RECT 115.85 291.47 116.01 293.06 ;
      RECT 115.13 292.38 116.01 292.54 ;
      RECT 115.85 294.86 116.01 296.45 ;
      RECT 115.13 295.38 116.01 295.54 ;
      RECT 115.85 298.27 116.01 299.86 ;
      RECT 115.13 299.18 116.01 299.34 ;
      RECT 115.85 301.66 116.01 303.25 ;
      RECT 115.13 302.18 116.01 302.34 ;
      RECT 115.85 305.07 116.01 306.66 ;
      RECT 115.13 305.98 116.01 306.14 ;
      RECT 115.85 308.46 116.01 310.05 ;
      RECT 115.13 308.98 116.01 309.14 ;
      RECT 115.85 311.87 116.01 313.46 ;
      RECT 115.13 312.78 116.01 312.94 ;
      RECT 115.85 315.26 116.01 316.85 ;
      RECT 115.13 315.78 116.01 315.94 ;
      RECT 115.85 318.67 116.01 320.26 ;
      RECT 115.13 319.58 116.01 319.74 ;
      RECT 115.85 322.06 116.01 323.65 ;
      RECT 115.13 322.58 116.01 322.74 ;
      RECT 115.85 325.47 116.01 327.06 ;
      RECT 115.13 326.38 116.01 326.54 ;
      RECT 115.85 328.86 116.01 330.45 ;
      RECT 115.13 329.38 116.01 329.54 ;
      RECT 115.85 332.27 116.01 333.86 ;
      RECT 115.13 333.18 116.01 333.34 ;
      RECT 115.85 335.66 116.01 337.25 ;
      RECT 115.13 336.18 116.01 336.34 ;
      RECT 115.85 339.07 116.01 340.66 ;
      RECT 115.13 339.98 116.01 340.14 ;
      RECT 115.85 342.46 116.01 344.05 ;
      RECT 115.13 342.98 116.01 343.14 ;
      RECT 115.85 345.87 116.01 347.46 ;
      RECT 115.13 346.78 116.01 346.94 ;
      RECT 115.85 349.26 116.01 350.85 ;
      RECT 115.13 349.78 116.01 349.94 ;
      RECT 115.85 352.67 116.01 354.26 ;
      RECT 115.13 353.58 116.01 353.74 ;
      RECT 115.85 356.06 116.01 357.65 ;
      RECT 115.13 356.58 116.01 356.74 ;
      RECT 115.85 359.47 116.01 361.06 ;
      RECT 115.13 360.38 116.01 360.54 ;
      RECT 115.85 362.86 116.01 364.45 ;
      RECT 115.13 363.38 116.01 363.54 ;
      RECT 115.85 366.27 116.01 367.86 ;
      RECT 115.13 367.18 116.01 367.34 ;
      RECT 115.85 369.66 116.01 371.25 ;
      RECT 115.13 370.18 116.01 370.34 ;
      RECT 115.85 373.07 116.01 374.66 ;
      RECT 115.13 373.98 116.01 374.14 ;
      RECT 115.85 376.46 116.01 378.05 ;
      RECT 115.13 376.98 116.01 377.14 ;
      RECT 115.85 379.87 116.01 381.46 ;
      RECT 115.13 380.78 116.01 380.94 ;
      RECT 115.85 383.26 116.01 384.85 ;
      RECT 115.13 383.78 116.01 383.94 ;
      RECT 115.85 386.67 116.01 388.26 ;
      RECT 115.13 387.58 116.01 387.74 ;
      RECT 115.85 390.06 116.01 391.65 ;
      RECT 115.13 390.58 116.01 390.74 ;
      RECT 115.85 393.47 116.01 395.06 ;
      RECT 115.13 394.38 116.01 394.54 ;
      RECT 115.85 396.86 116.01 398.45 ;
      RECT 115.13 397.38 116.01 397.54 ;
      RECT 115.85 400.27 116.01 401.86 ;
      RECT 115.13 401.18 116.01 401.34 ;
      RECT 115.85 403.66 116.01 405.25 ;
      RECT 115.13 404.18 116.01 404.34 ;
      RECT 115.85 407.07 116.01 408.66 ;
      RECT 115.13 407.98 116.01 408.14 ;
      RECT 115.85 410.46 116.01 412.05 ;
      RECT 115.13 410.98 116.01 411.14 ;
      RECT 115.85 413.87 116.01 415.46 ;
      RECT 115.13 414.78 116.01 414.94 ;
      RECT 115.85 417.26 116.01 418.85 ;
      RECT 115.13 417.78 116.01 417.94 ;
      RECT 115.85 420.67 116.01 422.26 ;
      RECT 115.13 421.58 116.01 421.74 ;
      RECT 115.85 424.06 116.01 425.65 ;
      RECT 115.13 424.58 116.01 424.74 ;
      RECT 115.85 427.47 116.01 429.06 ;
      RECT 115.13 428.38 116.01 428.54 ;
      RECT 115.85 430.86 116.01 432.45 ;
      RECT 115.13 431.38 116.01 431.54 ;
      RECT 115.85 434.27 116.01 435.86 ;
      RECT 115.13 435.18 116.01 435.34 ;
      RECT 115.85 437.66 116.01 439.25 ;
      RECT 115.13 438.18 116.01 438.34 ;
      RECT 115.85 441.07 116.01 442.66 ;
      RECT 115.13 441.98 116.01 442.14 ;
      RECT 115.85 444.46 116.01 446.05 ;
      RECT 115.13 444.98 116.01 445.14 ;
      RECT 115.85 447.87 116.01 449.46 ;
      RECT 115.13 448.78 116.01 448.94 ;
      RECT 115.85 451.26 116.01 452.85 ;
      RECT 115.13 451.78 116.01 451.94 ;
      RECT 115.85 454.67 116.01 456.26 ;
      RECT 115.13 455.58 116.01 455.74 ;
      RECT 115.85 458.06 116.01 459.65 ;
      RECT 115.13 458.58 116.01 458.74 ;
      RECT 115.85 461.47 116.01 463.06 ;
      RECT 115.13 462.38 116.01 462.54 ;
      RECT 115.85 464.86 116.01 466.45 ;
      RECT 115.13 465.38 116.01 465.54 ;
      RECT 115.85 468.27 116.01 469.86 ;
      RECT 115.13 469.18 116.01 469.34 ;
      RECT 115.85 471.66 116.01 473.25 ;
      RECT 115.13 472.18 116.01 472.34 ;
      RECT 115.85 475.07 116.01 476.66 ;
      RECT 115.13 475.98 116.01 476.14 ;
      RECT 115.85 478.46 116.01 480.05 ;
      RECT 115.13 478.98 116.01 479.14 ;
      RECT 115.85 481.87 116.01 483.46 ;
      RECT 115.13 482.78 116.01 482.94 ;
      RECT 115.85 485.26 116.01 486.85 ;
      RECT 115.13 485.78 116.01 485.94 ;
      RECT 115.85 488.67 116.01 490.26 ;
      RECT 115.13 489.58 116.01 489.74 ;
      RECT 115.85 492.06 116.01 493.65 ;
      RECT 115.13 492.58 116.01 492.74 ;
      RECT 115.85 495.47 116.01 497.06 ;
      RECT 115.13 496.38 116.01 496.54 ;
      RECT 115.85 498.86 116.01 500.45 ;
      RECT 115.13 499.38 116.01 499.54 ;
      RECT 115.85 502.27 116.01 503.86 ;
      RECT 115.13 503.18 116.01 503.34 ;
      RECT 115.15 49.6 115.31 51.7 ;
      RECT 115.15 49.6 115.75 49.76 ;
      RECT 115.59 32.06 115.75 49.76 ;
      RECT 114.93 45.9 115.75 46.06 ;
      RECT 114.93 36.23 115.75 36.39 ;
      RECT 115.15 32.06 115.75 32.22 ;
      RECT 115.15 30.54 115.31 32.22 ;
      RECT 113.65 21.06 113.81 26.28 ;
      RECT 114.61 24.37 114.77 25.98 ;
      RECT 113.65 24.37 114.97 24.53 ;
      RECT 114.81 23.67 114.97 24.53 ;
      RECT 114.61 23.67 114.97 23.83 ;
      RECT 114.61 21.7 114.77 23.83 ;
      RECT 113.59 21.06 115.47 21.22 ;
      RECT 113.59 60.83 115.47 60.99 ;
      RECT 113.65 55.81 113.81 60.99 ;
      RECT 114.61 58.22 114.77 60.35 ;
      RECT 114.61 58.22 114.97 58.38 ;
      RECT 114.81 57.25 114.97 58.38 ;
      RECT 113.65 57.25 114.97 57.41 ;
      RECT 114.61 56.13 114.77 57.41 ;
      RECT 113.25 25.79 113.49 26.07 ;
      RECT 113.33 21.94 113.49 26.07 ;
      RECT 113.21 21.94 113.49 22.18 ;
      RECT 113.27 15.28 113.43 22.18 ;
      RECT 115.19 15.28 115.35 20.88 ;
      RECT 114.23 15.28 114.39 20.88 ;
      RECT 113.27 17.14 115.35 17.3 ;
      RECT 113.27 35.91 115.35 36.07 ;
      RECT 115.19 32.85 115.35 36.07 ;
      RECT 114.23 27.43 114.39 36.07 ;
      RECT 113.27 32.85 113.43 36.07 ;
      RECT 114.23 27.43 115.29 27.59 ;
      RECT 115.13 23.41 115.29 27.59 ;
      RECT 114.13 26.14 115.29 26.3 ;
      RECT 115.09 25 115.29 26.3 ;
      RECT 114.13 25.01 114.29 26.3 ;
      RECT 114.13 21.38 114.29 23.81 ;
      RECT 115.09 21.38 115.25 23.55 ;
      RECT 114.13 21.38 115.25 21.54 ;
      RECT 114.13 60.51 115.25 60.67 ;
      RECT 115.09 58.5 115.25 60.67 ;
      RECT 115.13 55.81 115.25 60.67 ;
      RECT 114.13 58.24 114.29 60.67 ;
      RECT 115.15 54.64 115.29 58.64 ;
      RECT 115.09 55.81 115.31 57.09 ;
      RECT 115.15 54.64 115.31 57.09 ;
      RECT 114.13 55.81 114.29 57.09 ;
      RECT 114.13 55.81 115.31 55.97 ;
      RECT 114.23 54.64 115.31 54.8 ;
      RECT 114.23 46.22 114.39 54.8 ;
      RECT 115.19 46.22 115.35 49.44 ;
      RECT 113.27 46.22 113.43 49.44 ;
      RECT 113.27 46.22 115.35 46.38 ;
      RECT 115.19 61.17 115.35 66.77 ;
      RECT 114.23 61.17 114.39 66.77 ;
      RECT 113.27 59.87 113.43 66.77 ;
      RECT 113.27 64.75 115.35 64.91 ;
      RECT 113.21 59.87 113.49 60.11 ;
      RECT 113.33 56.02 113.49 60.11 ;
      RECT 113.25 56.02 113.49 56.3 ;
      RECT 114.23 10.09 114.39 14.2 ;
      RECT 114.23 12.9 115.29 13.06 ;
      RECT 115.13 12.19 115.29 13.06 ;
      RECT 115.11 41.08 115.27 45.17 ;
      RECT 114.95 41.08 115.27 41.24 ;
      RECT 114.71 14.52 114.87 16.86 ;
      RECT 114.84 13.22 115 14.84 ;
      RECT 114.71 31.09 114.87 35.75 ;
      RECT 114.71 32.25 114.97 32.53 ;
      RECT 112.93 26.46 114.95 26.62 ;
      RECT 112.93 25.35 113.09 26.62 ;
      RECT 113.01 22.91 113.17 25.51 ;
      RECT 113.01 56.46 113.17 59.14 ;
      RECT 112.93 55.49 113.09 56.62 ;
      RECT 112.93 55.49 114.95 55.65 ;
      RECT 114.71 49.75 114.91 51.3 ;
      RECT 114.71 46.54 114.87 51.3 ;
      RECT 113.59 55.09 114.85 55.25 ;
      RECT 113.59 49.77 113.75 55.25 ;
      RECT 112.87 49.77 113.75 49.93 ;
      RECT 112.87 32.48 113.03 49.93 ;
      RECT 112.87 45.9 113.69 46.06 ;
      RECT 112.87 36.23 113.69 36.39 ;
      RECT 112.87 32.48 113.75 32.64 ;
      RECT 113.59 27.04 113.75 32.64 ;
      RECT 113.59 27.04 114.85 27.2 ;
      RECT 113.97 45.9 114.77 46.06 ;
      RECT 114.61 44.89 114.77 46.06 ;
      RECT 114.63 38.57 114.79 45.17 ;
      RECT 113.83 38.57 113.99 45.17 ;
      RECT 113.83 38.57 114.29 38.73 ;
      RECT 114.13 36.23 114.29 38.73 ;
      RECT 113.97 36.23 114.65 36.39 ;
      RECT 113.75 32.85 113.91 35.75 ;
      RECT 113.91 31.09 114.07 33.01 ;
      RECT 113.91 49.44 114.07 51.3 ;
      RECT 113.75 46.54 113.91 49.6 ;
      RECT 113.33 12.8 113.99 13.06 ;
      RECT 113.33 12.19 113.57 13.06 ;
      RECT 113.75 14.52 113.91 16.86 ;
      RECT 113.62 13.22 113.78 14.84 ;
      RECT 113.35 41.08 113.51 45.17 ;
      RECT 113.35 41.08 113.67 41.24 ;
      RECT 112.53 17.6 112.69 23.81 ;
      RECT 112.05 22.38 113.17 22.54 ;
      RECT 112.53 58.24 112.69 64 ;
      RECT 112.05 59.51 113.17 59.67 ;
      RECT 112.95 27.37 113.11 31.49 ;
      RECT 112.11 27.37 112.27 31.49 ;
      RECT 112.11 27.37 113.11 27.53 ;
      RECT 112.53 24.64 112.69 27.53 ;
      RECT 112.53 54.16 112.69 57.42 ;
      RECT 112.11 54.16 113.11 54.88 ;
      RECT 112.95 50.8 113.11 54.88 ;
      RECT 112.11 50.8 112.27 54.88 ;
      RECT 110.37 55.09 111.63 55.25 ;
      RECT 111.47 49.77 111.63 55.25 ;
      RECT 111.47 49.77 112.35 49.93 ;
      RECT 112.19 32.48 112.35 49.93 ;
      RECT 111.53 45.9 112.35 46.06 ;
      RECT 111.53 36.23 112.35 36.39 ;
      RECT 111.47 32.48 112.35 32.64 ;
      RECT 111.47 27.04 111.63 32.64 ;
      RECT 110.37 27.04 111.63 27.2 ;
      RECT 110.27 26.46 112.29 26.62 ;
      RECT 112.13 25.35 112.29 26.62 ;
      RECT 112.05 22.91 112.21 25.51 ;
      RECT 112.05 56.46 112.21 59.14 ;
      RECT 112.13 55.49 112.29 56.62 ;
      RECT 110.27 55.49 112.29 55.65 ;
      RECT 111.64 9.18 111.8 14.23 ;
      RECT 110.11 9.18 110.27 14.23 ;
      RECT 110.11 11.85 111.8 12.01 ;
      RECT 110.11 9.18 111.8 9.34 ;
      RECT 110.58 7.64 111.26 9.34 ;
      RECT 109.85 7.64 112.13 8.28 ;
      RECT 111.73 25.79 111.97 26.07 ;
      RECT 111.73 21.94 111.89 26.07 ;
      RECT 111.73 21.94 112.01 22.18 ;
      RECT 111.79 15.28 111.95 22.18 ;
      RECT 110.83 15.28 110.99 20.88 ;
      RECT 109.87 15.28 110.03 20.88 ;
      RECT 109.87 17.14 111.95 17.3 ;
      RECT 111.79 59.87 111.95 66.77 ;
      RECT 110.83 61.17 110.99 66.77 ;
      RECT 109.87 61.17 110.03 66.77 ;
      RECT 109.87 64.75 111.95 64.91 ;
      RECT 111.73 59.87 112.01 60.11 ;
      RECT 111.73 56.02 111.89 60.11 ;
      RECT 111.73 56.02 111.97 56.3 ;
      RECT 109.87 35.91 111.95 36.07 ;
      RECT 111.79 32.85 111.95 36.07 ;
      RECT 110.83 27.43 110.99 36.07 ;
      RECT 109.87 32.85 110.03 36.07 ;
      RECT 109.93 27.43 110.99 27.59 ;
      RECT 109.93 23.41 110.09 27.59 ;
      RECT 109.93 26.14 111.09 26.3 ;
      RECT 110.93 25.01 111.09 26.3 ;
      RECT 109.93 25 110.13 26.3 ;
      RECT 110.93 21.38 111.09 23.81 ;
      RECT 109.97 21.38 110.13 23.55 ;
      RECT 109.97 21.38 111.09 21.54 ;
      RECT 109.97 60.51 111.09 60.67 ;
      RECT 110.93 58.24 111.09 60.67 ;
      RECT 109.97 58.5 110.13 60.67 ;
      RECT 109.93 55.81 110.09 58.64 ;
      RECT 110.93 55.81 111.09 57.09 ;
      RECT 109.91 55.81 110.13 57.09 ;
      RECT 109.91 55.81 111.09 55.97 ;
      RECT 109.91 54.64 110.07 57.09 ;
      RECT 109.91 54.64 110.99 54.8 ;
      RECT 110.83 46.22 110.99 54.8 ;
      RECT 111.79 46.22 111.95 49.44 ;
      RECT 109.87 46.22 110.03 49.44 ;
      RECT 109.87 46.22 111.95 46.38 ;
      RECT 111.71 41.08 111.87 45.17 ;
      RECT 111.55 41.08 111.87 41.24 ;
      RECT 111.41 21.06 111.57 26.28 ;
      RECT 110.45 24.37 110.61 25.98 ;
      RECT 110.25 24.37 111.57 24.53 ;
      RECT 110.25 23.67 110.41 24.53 ;
      RECT 110.25 23.67 110.61 23.83 ;
      RECT 110.45 21.7 110.61 23.83 ;
      RECT 109.75 21.06 111.63 21.22 ;
      RECT 109.75 60.83 111.63 60.99 ;
      RECT 111.41 55.81 111.57 60.99 ;
      RECT 110.45 58.22 110.61 60.35 ;
      RECT 110.25 58.22 110.61 58.38 ;
      RECT 110.25 57.25 110.41 58.38 ;
      RECT 110.25 57.25 111.57 57.41 ;
      RECT 110.45 56.13 110.61 57.41 ;
      RECT 111.31 32.85 111.47 35.75 ;
      RECT 111.15 31.09 111.31 33.01 ;
      RECT 111.15 49.44 111.31 51.3 ;
      RECT 111.31 46.54 111.47 49.6 ;
      RECT 111.23 38.57 111.39 45.17 ;
      RECT 110.93 38.57 111.39 38.73 ;
      RECT 110.93 36.23 111.09 38.73 ;
      RECT 110.57 36.23 111.25 36.39 ;
      RECT 110.45 45.9 111.25 46.06 ;
      RECT 110.45 44.89 110.61 46.06 ;
      RECT 110.43 38.57 110.59 45.17 ;
      RECT 110.35 31.09 110.51 35.75 ;
      RECT 110.25 32.25 110.51 32.53 ;
      RECT 110.31 49.75 110.51 51.3 ;
      RECT 110.35 46.54 110.51 51.3 ;
      RECT 109.38 70.94 110.3 71.18 ;
      RECT 96.66 70.96 110.3 71.16 ;
      RECT 108.21 74.7 108.81 75.05 ;
      RECT 109.38 74.74 110.3 74.98 ;
      RECT 108.21 74.76 110.3 74.96 ;
      RECT 108.21 77.67 108.81 78.02 ;
      RECT 109.38 77.74 110.3 77.98 ;
      RECT 108.21 77.76 110.3 77.96 ;
      RECT 108.21 81.5 108.81 81.85 ;
      RECT 109.38 81.54 110.3 81.78 ;
      RECT 108.21 81.56 110.3 81.76 ;
      RECT 108.3 84.43 108.81 84.83 ;
      RECT 109.38 84.54 110.3 84.78 ;
      RECT 96.66 84.56 110.3 84.76 ;
      RECT 108.21 88.3 108.81 88.65 ;
      RECT 109.38 88.34 110.3 88.58 ;
      RECT 108.21 88.36 110.3 88.56 ;
      RECT 108.21 91.27 108.81 91.62 ;
      RECT 109.38 91.34 110.3 91.58 ;
      RECT 108.21 91.36 110.3 91.56 ;
      RECT 108.21 95.1 108.81 95.45 ;
      RECT 109.38 95.14 110.3 95.38 ;
      RECT 108.21 95.16 110.3 95.36 ;
      RECT 108.3 98.03 108.81 98.43 ;
      RECT 109.38 98.14 110.3 98.38 ;
      RECT 96.66 98.16 110.3 98.36 ;
      RECT 108.21 101.9 108.81 102.25 ;
      RECT 109.38 101.94 110.3 102.18 ;
      RECT 108.21 101.96 110.3 102.16 ;
      RECT 108.21 104.87 108.81 105.22 ;
      RECT 109.38 104.94 110.3 105.18 ;
      RECT 108.21 104.96 110.3 105.16 ;
      RECT 108.21 108.7 108.81 109.05 ;
      RECT 109.38 108.74 110.3 108.98 ;
      RECT 108.21 108.76 110.3 108.96 ;
      RECT 108.3 111.63 108.81 112.03 ;
      RECT 109.38 111.74 110.3 111.98 ;
      RECT 96.66 111.76 110.3 111.96 ;
      RECT 108.21 115.5 108.81 115.85 ;
      RECT 109.38 115.54 110.3 115.78 ;
      RECT 108.21 115.56 110.3 115.76 ;
      RECT 108.21 118.47 108.81 118.82 ;
      RECT 109.38 118.54 110.3 118.78 ;
      RECT 108.21 118.56 110.3 118.76 ;
      RECT 108.21 122.3 108.81 122.65 ;
      RECT 109.38 122.34 110.3 122.58 ;
      RECT 108.21 122.36 110.3 122.56 ;
      RECT 108.3 125.23 108.81 125.63 ;
      RECT 109.38 125.34 110.3 125.58 ;
      RECT 96.66 125.36 110.3 125.56 ;
      RECT 108.21 129.1 108.81 129.45 ;
      RECT 109.38 129.14 110.3 129.38 ;
      RECT 108.21 129.16 110.3 129.36 ;
      RECT 108.21 132.07 108.81 132.42 ;
      RECT 109.38 132.14 110.3 132.38 ;
      RECT 108.21 132.16 110.3 132.36 ;
      RECT 108.21 135.9 108.81 136.25 ;
      RECT 109.38 135.94 110.3 136.18 ;
      RECT 108.21 135.96 110.3 136.16 ;
      RECT 108.3 138.83 108.81 139.23 ;
      RECT 109.38 138.94 110.3 139.18 ;
      RECT 96.66 138.96 110.3 139.16 ;
      RECT 108.21 142.7 108.81 143.05 ;
      RECT 109.38 142.74 110.3 142.98 ;
      RECT 108.21 142.76 110.3 142.96 ;
      RECT 108.21 145.67 108.81 146.02 ;
      RECT 109.38 145.74 110.3 145.98 ;
      RECT 108.21 145.76 110.3 145.96 ;
      RECT 108.21 149.5 108.81 149.85 ;
      RECT 109.38 149.54 110.3 149.78 ;
      RECT 108.21 149.56 110.3 149.76 ;
      RECT 108.3 152.43 108.81 152.83 ;
      RECT 109.38 152.54 110.3 152.78 ;
      RECT 96.66 152.56 110.3 152.76 ;
      RECT 108.21 156.3 108.81 156.65 ;
      RECT 109.38 156.34 110.3 156.58 ;
      RECT 108.21 156.36 110.3 156.56 ;
      RECT 108.21 159.27 108.81 159.62 ;
      RECT 109.38 159.34 110.3 159.58 ;
      RECT 108.21 159.36 110.3 159.56 ;
      RECT 108.21 163.1 108.81 163.45 ;
      RECT 109.38 163.14 110.3 163.38 ;
      RECT 108.21 163.16 110.3 163.36 ;
      RECT 108.3 166.03 108.81 166.43 ;
      RECT 109.38 166.14 110.3 166.38 ;
      RECT 96.66 166.16 110.3 166.36 ;
      RECT 108.21 169.9 108.81 170.25 ;
      RECT 109.38 169.94 110.3 170.18 ;
      RECT 108.21 169.96 110.3 170.16 ;
      RECT 108.21 172.87 108.81 173.22 ;
      RECT 109.38 172.94 110.3 173.18 ;
      RECT 108.21 172.96 110.3 173.16 ;
      RECT 108.21 176.7 108.81 177.05 ;
      RECT 109.38 176.74 110.3 176.98 ;
      RECT 108.21 176.76 110.3 176.96 ;
      RECT 108.32 179.65 108.7 180.04 ;
      RECT 109.38 179.74 110.3 179.98 ;
      RECT 96.66 179.76 110.3 179.96 ;
      RECT 108.21 183.5 108.81 183.85 ;
      RECT 109.38 183.54 110.3 183.78 ;
      RECT 108.21 183.56 110.3 183.76 ;
      RECT 108.21 186.47 108.81 186.82 ;
      RECT 109.38 186.54 110.3 186.78 ;
      RECT 108.21 186.56 110.3 186.76 ;
      RECT 108.21 190.3 108.81 190.65 ;
      RECT 109.38 190.34 110.3 190.58 ;
      RECT 108.21 190.36 110.3 190.56 ;
      RECT 108.3 193.23 108.81 193.63 ;
      RECT 109.38 193.34 110.3 193.58 ;
      RECT 96.66 193.36 110.3 193.56 ;
      RECT 108.21 197.1 108.81 197.45 ;
      RECT 109.38 197.14 110.3 197.38 ;
      RECT 108.21 197.16 110.3 197.36 ;
      RECT 108.21 200.07 108.81 200.42 ;
      RECT 109.38 200.14 110.3 200.38 ;
      RECT 108.21 200.16 110.3 200.36 ;
      RECT 108.21 203.9 108.81 204.25 ;
      RECT 109.38 203.94 110.3 204.18 ;
      RECT 108.21 203.96 110.3 204.16 ;
      RECT 108.3 206.83 108.81 207.23 ;
      RECT 109.38 206.94 110.3 207.18 ;
      RECT 96.66 206.96 110.3 207.16 ;
      RECT 108.21 210.7 108.81 211.05 ;
      RECT 109.38 210.74 110.3 210.98 ;
      RECT 108.21 210.76 110.3 210.96 ;
      RECT 108.21 213.67 108.81 214.02 ;
      RECT 109.38 213.74 110.3 213.98 ;
      RECT 108.21 213.76 110.3 213.96 ;
      RECT 108.21 217.5 108.81 217.85 ;
      RECT 109.38 217.54 110.3 217.78 ;
      RECT 108.21 217.56 110.3 217.76 ;
      RECT 108.3 220.43 108.81 220.83 ;
      RECT 109.38 220.54 110.3 220.78 ;
      RECT 96.66 220.56 110.3 220.76 ;
      RECT 108.21 224.3 108.81 224.65 ;
      RECT 109.38 224.34 110.3 224.58 ;
      RECT 108.21 224.36 110.3 224.56 ;
      RECT 108.21 227.27 108.81 227.62 ;
      RECT 109.38 227.34 110.3 227.58 ;
      RECT 108.21 227.36 110.3 227.56 ;
      RECT 108.21 231.1 108.81 231.45 ;
      RECT 109.38 231.14 110.3 231.38 ;
      RECT 108.21 231.16 110.3 231.36 ;
      RECT 108.3 234.03 108.81 234.43 ;
      RECT 109.38 234.14 110.3 234.38 ;
      RECT 96.66 234.16 110.3 234.36 ;
      RECT 108.21 237.9 108.81 238.25 ;
      RECT 109.38 237.94 110.3 238.18 ;
      RECT 108.21 237.96 110.3 238.16 ;
      RECT 108.21 240.87 108.81 241.22 ;
      RECT 109.38 240.94 110.3 241.18 ;
      RECT 108.21 240.96 110.3 241.16 ;
      RECT 108.21 244.7 108.81 245.05 ;
      RECT 109.38 244.74 110.3 244.98 ;
      RECT 108.21 244.76 110.3 244.96 ;
      RECT 108.3 247.63 108.81 248.03 ;
      RECT 109.38 247.74 110.3 247.98 ;
      RECT 96.66 247.76 110.3 247.96 ;
      RECT 108.21 251.5 108.81 251.85 ;
      RECT 109.38 251.54 110.3 251.78 ;
      RECT 108.21 251.56 110.3 251.76 ;
      RECT 108.21 254.47 108.81 254.82 ;
      RECT 109.38 254.54 110.3 254.78 ;
      RECT 108.21 254.56 110.3 254.76 ;
      RECT 108.21 258.3 108.81 258.65 ;
      RECT 109.38 258.34 110.3 258.58 ;
      RECT 108.21 258.36 110.3 258.56 ;
      RECT 108.3 261.23 108.81 261.63 ;
      RECT 109.38 261.34 110.3 261.58 ;
      RECT 96.66 261.36 110.3 261.56 ;
      RECT 108.21 265.1 108.81 265.45 ;
      RECT 109.38 265.14 110.3 265.38 ;
      RECT 108.21 265.16 110.3 265.36 ;
      RECT 108.21 268.07 108.81 268.42 ;
      RECT 109.38 268.14 110.3 268.38 ;
      RECT 108.21 268.16 110.3 268.36 ;
      RECT 108.21 271.9 108.81 272.25 ;
      RECT 109.38 271.94 110.3 272.18 ;
      RECT 108.21 271.96 110.3 272.16 ;
      RECT 108.3 274.83 108.81 275.23 ;
      RECT 109.38 274.94 110.3 275.18 ;
      RECT 96.66 274.96 110.3 275.16 ;
      RECT 108.21 278.7 108.81 279.05 ;
      RECT 109.38 278.74 110.3 278.98 ;
      RECT 108.21 278.76 110.3 278.96 ;
      RECT 108.21 281.67 108.81 282.02 ;
      RECT 109.38 281.74 110.3 281.98 ;
      RECT 108.21 281.76 110.3 281.96 ;
      RECT 108.21 285.5 108.81 285.85 ;
      RECT 109.38 285.54 110.3 285.78 ;
      RECT 108.21 285.56 110.3 285.76 ;
      RECT 108.32 288.45 108.7 288.84 ;
      RECT 109.38 288.54 110.3 288.78 ;
      RECT 96.66 288.56 110.3 288.76 ;
      RECT 108.21 292.3 108.81 292.65 ;
      RECT 109.38 292.34 110.3 292.58 ;
      RECT 108.21 292.36 110.3 292.56 ;
      RECT 108.21 295.27 108.81 295.62 ;
      RECT 109.38 295.34 110.3 295.58 ;
      RECT 108.21 295.36 110.3 295.56 ;
      RECT 108.21 299.1 108.81 299.45 ;
      RECT 109.38 299.14 110.3 299.38 ;
      RECT 108.21 299.16 110.3 299.36 ;
      RECT 108.3 302.03 108.81 302.43 ;
      RECT 109.38 302.14 110.3 302.38 ;
      RECT 96.66 302.16 110.3 302.36 ;
      RECT 108.21 305.9 108.81 306.25 ;
      RECT 109.38 305.94 110.3 306.18 ;
      RECT 108.21 305.96 110.3 306.16 ;
      RECT 108.21 308.87 108.81 309.22 ;
      RECT 109.38 308.94 110.3 309.18 ;
      RECT 108.21 308.96 110.3 309.16 ;
      RECT 108.21 312.7 108.81 313.05 ;
      RECT 109.38 312.74 110.3 312.98 ;
      RECT 108.21 312.76 110.3 312.96 ;
      RECT 108.3 315.63 108.81 316.03 ;
      RECT 109.38 315.74 110.3 315.98 ;
      RECT 96.66 315.76 110.3 315.96 ;
      RECT 108.21 319.5 108.81 319.85 ;
      RECT 109.38 319.54 110.3 319.78 ;
      RECT 108.21 319.56 110.3 319.76 ;
      RECT 108.21 322.47 108.81 322.82 ;
      RECT 109.38 322.54 110.3 322.78 ;
      RECT 108.21 322.56 110.3 322.76 ;
      RECT 108.21 326.3 108.81 326.65 ;
      RECT 109.38 326.34 110.3 326.58 ;
      RECT 108.21 326.36 110.3 326.56 ;
      RECT 108.3 329.23 108.81 329.63 ;
      RECT 109.38 329.34 110.3 329.58 ;
      RECT 96.66 329.36 110.3 329.56 ;
      RECT 108.21 333.1 108.81 333.45 ;
      RECT 109.38 333.14 110.3 333.38 ;
      RECT 108.21 333.16 110.3 333.36 ;
      RECT 108.21 336.07 108.81 336.42 ;
      RECT 109.38 336.14 110.3 336.38 ;
      RECT 108.21 336.16 110.3 336.36 ;
      RECT 108.21 339.9 108.81 340.25 ;
      RECT 109.38 339.94 110.3 340.18 ;
      RECT 108.21 339.96 110.3 340.16 ;
      RECT 108.3 342.83 108.81 343.23 ;
      RECT 109.38 342.94 110.3 343.18 ;
      RECT 96.66 342.96 110.3 343.16 ;
      RECT 108.21 346.7 108.81 347.05 ;
      RECT 109.38 346.74 110.3 346.98 ;
      RECT 108.21 346.76 110.3 346.96 ;
      RECT 108.21 349.67 108.81 350.02 ;
      RECT 109.38 349.74 110.3 349.98 ;
      RECT 108.21 349.76 110.3 349.96 ;
      RECT 108.21 353.5 108.81 353.85 ;
      RECT 109.38 353.54 110.3 353.78 ;
      RECT 108.21 353.56 110.3 353.76 ;
      RECT 108.3 356.43 108.81 356.83 ;
      RECT 109.38 356.54 110.3 356.78 ;
      RECT 96.66 356.56 110.3 356.76 ;
      RECT 108.21 360.3 108.81 360.65 ;
      RECT 109.38 360.34 110.3 360.58 ;
      RECT 108.21 360.36 110.3 360.56 ;
      RECT 108.21 363.27 108.81 363.62 ;
      RECT 109.38 363.34 110.3 363.58 ;
      RECT 108.21 363.36 110.3 363.56 ;
      RECT 108.21 367.1 108.81 367.45 ;
      RECT 109.38 367.14 110.3 367.38 ;
      RECT 108.21 367.16 110.3 367.36 ;
      RECT 108.3 370.03 108.81 370.43 ;
      RECT 109.38 370.14 110.3 370.38 ;
      RECT 96.66 370.16 110.3 370.36 ;
      RECT 108.21 373.9 108.81 374.25 ;
      RECT 109.38 373.94 110.3 374.18 ;
      RECT 108.21 373.96 110.3 374.16 ;
      RECT 108.21 376.87 108.81 377.22 ;
      RECT 109.38 376.94 110.3 377.18 ;
      RECT 108.21 376.96 110.3 377.16 ;
      RECT 108.21 380.7 108.81 381.05 ;
      RECT 109.38 380.74 110.3 380.98 ;
      RECT 108.21 380.76 110.3 380.96 ;
      RECT 108.3 383.63 108.81 384.03 ;
      RECT 109.38 383.74 110.3 383.98 ;
      RECT 96.66 383.76 110.3 383.96 ;
      RECT 108.21 387.5 108.81 387.85 ;
      RECT 109.38 387.54 110.3 387.78 ;
      RECT 108.21 387.56 110.3 387.76 ;
      RECT 108.21 390.47 108.81 390.82 ;
      RECT 109.38 390.54 110.3 390.78 ;
      RECT 108.21 390.56 110.3 390.76 ;
      RECT 108.21 394.3 108.81 394.65 ;
      RECT 109.38 394.34 110.3 394.58 ;
      RECT 108.21 394.36 110.3 394.56 ;
      RECT 108.32 397.25 108.7 397.64 ;
      RECT 109.38 397.34 110.3 397.58 ;
      RECT 96.66 397.36 110.3 397.56 ;
      RECT 108.21 401.1 108.81 401.45 ;
      RECT 109.38 401.14 110.3 401.38 ;
      RECT 108.21 401.16 110.3 401.36 ;
      RECT 108.21 404.07 108.81 404.42 ;
      RECT 109.38 404.14 110.3 404.38 ;
      RECT 108.21 404.16 110.3 404.36 ;
      RECT 108.21 407.9 108.81 408.25 ;
      RECT 109.38 407.94 110.3 408.18 ;
      RECT 108.21 407.96 110.3 408.16 ;
      RECT 108.3 410.83 108.81 411.23 ;
      RECT 109.38 410.94 110.3 411.18 ;
      RECT 96.66 410.96 110.3 411.16 ;
      RECT 108.21 414.7 108.81 415.05 ;
      RECT 109.38 414.74 110.3 414.98 ;
      RECT 108.21 414.76 110.3 414.96 ;
      RECT 108.21 417.67 108.81 418.02 ;
      RECT 109.38 417.74 110.3 417.98 ;
      RECT 108.21 417.76 110.3 417.96 ;
      RECT 108.21 421.5 108.81 421.85 ;
      RECT 109.38 421.54 110.3 421.78 ;
      RECT 108.21 421.56 110.3 421.76 ;
      RECT 108.3 424.43 108.81 424.83 ;
      RECT 109.38 424.54 110.3 424.78 ;
      RECT 96.66 424.56 110.3 424.76 ;
      RECT 108.21 428.3 108.81 428.65 ;
      RECT 109.38 428.34 110.3 428.58 ;
      RECT 108.21 428.36 110.3 428.56 ;
      RECT 108.21 431.27 108.81 431.62 ;
      RECT 109.38 431.34 110.3 431.58 ;
      RECT 108.21 431.36 110.3 431.56 ;
      RECT 108.21 435.1 108.81 435.45 ;
      RECT 109.38 435.14 110.3 435.38 ;
      RECT 108.21 435.16 110.3 435.36 ;
      RECT 108.3 438.03 108.81 438.43 ;
      RECT 109.38 438.14 110.3 438.38 ;
      RECT 96.66 438.16 110.3 438.36 ;
      RECT 108.21 441.9 108.81 442.25 ;
      RECT 109.38 441.94 110.3 442.18 ;
      RECT 108.21 441.96 110.3 442.16 ;
      RECT 108.21 444.87 108.81 445.22 ;
      RECT 109.38 444.94 110.3 445.18 ;
      RECT 108.21 444.96 110.3 445.16 ;
      RECT 108.21 448.7 108.81 449.05 ;
      RECT 109.38 448.74 110.3 448.98 ;
      RECT 108.21 448.76 110.3 448.96 ;
      RECT 108.3 451.63 108.81 452.03 ;
      RECT 109.38 451.74 110.3 451.98 ;
      RECT 96.66 451.76 110.3 451.96 ;
      RECT 108.21 455.5 108.81 455.85 ;
      RECT 109.38 455.54 110.3 455.78 ;
      RECT 108.21 455.56 110.3 455.76 ;
      RECT 108.21 458.47 108.81 458.82 ;
      RECT 109.38 458.54 110.3 458.78 ;
      RECT 108.21 458.56 110.3 458.76 ;
      RECT 108.21 462.3 108.81 462.65 ;
      RECT 109.38 462.34 110.3 462.58 ;
      RECT 108.21 462.36 110.3 462.56 ;
      RECT 108.3 465.23 108.81 465.63 ;
      RECT 109.38 465.34 110.3 465.58 ;
      RECT 96.66 465.36 110.3 465.56 ;
      RECT 108.21 469.1 108.81 469.45 ;
      RECT 109.38 469.14 110.3 469.38 ;
      RECT 108.21 469.16 110.3 469.36 ;
      RECT 108.21 472.07 108.81 472.42 ;
      RECT 109.38 472.14 110.3 472.38 ;
      RECT 108.21 472.16 110.3 472.36 ;
      RECT 108.21 475.9 108.81 476.25 ;
      RECT 109.38 475.94 110.3 476.18 ;
      RECT 108.21 475.96 110.3 476.16 ;
      RECT 108.3 478.83 108.81 479.23 ;
      RECT 109.38 478.94 110.3 479.18 ;
      RECT 96.66 478.96 110.3 479.16 ;
      RECT 108.21 482.7 108.81 483.05 ;
      RECT 109.38 482.74 110.3 482.98 ;
      RECT 108.21 482.76 110.3 482.96 ;
      RECT 108.21 485.67 108.81 486.02 ;
      RECT 109.38 485.74 110.3 485.98 ;
      RECT 108.21 485.76 110.3 485.96 ;
      RECT 108.21 489.5 108.81 489.85 ;
      RECT 109.38 489.54 110.3 489.78 ;
      RECT 108.21 489.56 110.3 489.76 ;
      RECT 108.3 492.43 108.81 492.83 ;
      RECT 109.38 492.54 110.3 492.78 ;
      RECT 96.66 492.56 110.3 492.76 ;
      RECT 108.21 496.3 108.81 496.65 ;
      RECT 109.38 496.34 110.3 496.58 ;
      RECT 108.21 496.36 110.3 496.56 ;
      RECT 108.21 499.27 108.81 499.62 ;
      RECT 109.38 499.34 110.3 499.58 ;
      RECT 108.21 499.36 110.3 499.56 ;
      RECT 108.21 503.1 108.81 503.45 ;
      RECT 109.38 503.14 110.3 503.38 ;
      RECT 108.21 503.16 110.3 503.36 ;
      RECT 109.91 49.6 110.07 51.7 ;
      RECT 109.47 49.6 110.07 49.76 ;
      RECT 109.47 32.06 109.63 49.76 ;
      RECT 109.47 45.9 110.29 46.06 ;
      RECT 109.47 36.23 110.29 36.39 ;
      RECT 109.47 32.06 110.07 32.22 ;
      RECT 109.91 30.54 110.07 32.22 ;
      RECT 109.95 41.08 110.11 45.17 ;
      RECT 109.95 41.08 110.27 41.24 ;
      RECT 109.13 31.49 109.29 32.02 ;
      RECT 108.67 31.49 109.75 31.65 ;
      RECT 109.59 27.38 109.75 31.65 ;
      RECT 108.67 27.38 108.83 31.65 ;
      RECT 108.67 27.38 109.75 27.54 ;
      RECT 109.13 26.91 109.29 27.54 ;
      RECT 108.67 51.06 109.75 55.29 ;
      RECT 109.13 50.27 109.29 55.29 ;
      RECT 109.49 49.92 109.65 50.9 ;
      RECT 108.77 49.92 108.93 50.9 ;
      RECT 108.77 49.92 109.65 50.08 ;
      RECT 109.13 45.65 109.29 50.08 ;
      RECT 107.87 12.34 108.15 12.62 ;
      RECT 106.95 12.34 107.23 12.62 ;
      RECT 104.39 12.34 104.67 12.62 ;
      RECT 103.47 12.34 103.75 12.62 ;
      RECT 101.07 12.34 101.35 12.62 ;
      RECT 100.15 12.34 100.43 12.62 ;
      RECT 107.99 11.75 108.15 12.62 ;
      RECT 106.95 11.75 107.11 12.62 ;
      RECT 104.51 11.75 104.67 12.62 ;
      RECT 103.47 11.75 103.63 12.62 ;
      RECT 101.19 11.75 101.35 12.62 ;
      RECT 100.15 11.75 100.31 12.62 ;
      RECT 109.13 8.38 109.29 12.03 ;
      RECT 108.03 9.02 108.19 12.03 ;
      RECT 106.83 9.02 106.99 12.03 ;
      RECT 105.73 8.38 105.89 12.03 ;
      RECT 104.63 9.02 104.79 12.03 ;
      RECT 103.43 9.02 103.59 12.03 ;
      RECT 102.33 8.38 102.49 12.03 ;
      RECT 101.23 9.02 101.39 12.03 ;
      RECT 100.03 9.02 100.19 12.03 ;
      RECT 98.93 8.38 99.09 12.03 ;
      RECT 98.93 9.02 109.29 9.3 ;
      RECT 108.45 8.38 108.69 9.3 ;
      RECT 107.77 8.38 108.01 9.3 ;
      RECT 107.02 8.38 107.26 9.3 ;
      RECT 106.33 8.38 106.57 9.3 ;
      RECT 105.05 8.38 105.29 9.3 ;
      RECT 104.36 8.38 104.6 9.3 ;
      RECT 103.61 8.38 103.85 9.3 ;
      RECT 102.93 8.38 103.17 9.3 ;
      RECT 101.65 8.38 101.89 9.3 ;
      RECT 100.97 8.38 101.21 9.3 ;
      RECT 100.22 8.38 100.46 9.3 ;
      RECT 99.53 8.38 99.77 9.3 ;
      RECT 108.35 49.6 108.51 51.7 ;
      RECT 108.35 49.6 108.95 49.76 ;
      RECT 108.79 32.06 108.95 49.76 ;
      RECT 108.13 45.9 108.95 46.06 ;
      RECT 108.13 36.23 108.95 36.39 ;
      RECT 108.35 32.06 108.95 32.22 ;
      RECT 108.35 30.54 108.51 32.22 ;
      RECT 106.85 21.06 107.01 26.28 ;
      RECT 107.81 24.37 107.97 25.98 ;
      RECT 106.85 24.37 108.17 24.53 ;
      RECT 108.01 23.67 108.17 24.53 ;
      RECT 107.81 23.67 108.17 23.83 ;
      RECT 107.81 21.7 107.97 23.83 ;
      RECT 106.79 21.06 108.67 21.22 ;
      RECT 106.79 60.83 108.67 60.99 ;
      RECT 106.85 55.81 107.01 60.99 ;
      RECT 107.81 58.22 107.97 60.35 ;
      RECT 107.81 58.22 108.17 58.38 ;
      RECT 108.01 57.25 108.17 58.38 ;
      RECT 106.85 57.25 108.17 57.41 ;
      RECT 107.81 56.13 107.97 57.41 ;
      RECT 106.45 25.79 106.69 26.07 ;
      RECT 106.53 21.94 106.69 26.07 ;
      RECT 106.41 21.94 106.69 22.18 ;
      RECT 106.47 15.28 106.63 22.18 ;
      RECT 108.39 15.28 108.55 20.88 ;
      RECT 107.43 15.28 107.59 20.88 ;
      RECT 106.47 17.14 108.55 17.3 ;
      RECT 106.47 35.91 108.55 36.07 ;
      RECT 108.39 32.85 108.55 36.07 ;
      RECT 107.43 27.43 107.59 36.07 ;
      RECT 106.47 32.85 106.63 36.07 ;
      RECT 107.43 27.43 108.49 27.59 ;
      RECT 108.33 23.41 108.49 27.59 ;
      RECT 107.33 26.14 108.49 26.3 ;
      RECT 108.29 25 108.49 26.3 ;
      RECT 107.33 25.01 107.49 26.3 ;
      RECT 107.33 21.38 107.49 23.81 ;
      RECT 108.29 21.38 108.45 23.55 ;
      RECT 107.33 21.38 108.45 21.54 ;
      RECT 107.33 60.51 108.45 60.67 ;
      RECT 108.29 58.5 108.45 60.67 ;
      RECT 108.33 55.81 108.45 60.67 ;
      RECT 107.33 58.24 107.49 60.67 ;
      RECT 108.35 54.64 108.49 58.64 ;
      RECT 108.29 55.81 108.51 57.09 ;
      RECT 108.35 54.64 108.51 57.09 ;
      RECT 107.33 55.81 107.49 57.09 ;
      RECT 107.33 55.81 108.51 55.97 ;
      RECT 107.43 54.64 108.51 54.8 ;
      RECT 107.43 46.22 107.59 54.8 ;
      RECT 108.39 46.22 108.55 49.44 ;
      RECT 106.47 46.22 106.63 49.44 ;
      RECT 106.47 46.22 108.55 46.38 ;
      RECT 108.39 61.17 108.55 66.77 ;
      RECT 107.43 61.17 107.59 66.77 ;
      RECT 106.47 59.87 106.63 66.77 ;
      RECT 106.47 64.75 108.55 64.91 ;
      RECT 106.41 59.87 106.69 60.11 ;
      RECT 106.53 56.02 106.69 60.11 ;
      RECT 106.45 56.02 106.69 56.3 ;
      RECT 107.43 10.09 107.59 14.2 ;
      RECT 107.43 12.9 108.49 13.06 ;
      RECT 108.33 12.19 108.49 13.06 ;
      RECT 108.31 41.08 108.47 45.17 ;
      RECT 108.15 41.08 108.47 41.24 ;
      RECT 107.91 14.52 108.07 16.86 ;
      RECT 108.04 13.22 108.2 14.84 ;
      RECT 107.91 31.09 108.07 35.75 ;
      RECT 107.91 32.25 108.17 32.53 ;
      RECT 106.13 26.46 108.15 26.62 ;
      RECT 106.13 25.35 106.29 26.62 ;
      RECT 106.21 22.91 106.37 25.51 ;
      RECT 106.21 56.46 106.37 59.14 ;
      RECT 106.13 55.49 106.29 56.62 ;
      RECT 106.13 55.49 108.15 55.65 ;
      RECT 107.91 49.75 108.11 51.3 ;
      RECT 107.91 46.54 108.07 51.3 ;
      RECT 106.79 55.09 108.05 55.25 ;
      RECT 106.79 49.77 106.95 55.25 ;
      RECT 106.07 49.77 106.95 49.93 ;
      RECT 106.07 32.48 106.23 49.93 ;
      RECT 106.07 45.9 106.89 46.06 ;
      RECT 106.07 36.23 106.89 36.39 ;
      RECT 106.07 32.48 106.95 32.64 ;
      RECT 106.79 27.04 106.95 32.64 ;
      RECT 106.79 27.04 108.05 27.2 ;
      RECT 107.17 45.9 107.97 46.06 ;
      RECT 107.81 44.89 107.97 46.06 ;
      RECT 107.83 38.57 107.99 45.17 ;
      RECT 107.03 38.57 107.19 45.17 ;
      RECT 107.03 38.57 107.49 38.73 ;
      RECT 107.33 36.23 107.49 38.73 ;
      RECT 107.17 36.23 107.85 36.39 ;
      RECT 106.95 32.85 107.11 35.75 ;
      RECT 107.11 31.09 107.27 33.01 ;
      RECT 107.11 49.44 107.27 51.3 ;
      RECT 106.95 46.54 107.11 49.6 ;
      RECT 106.53 12.8 107.19 13.06 ;
      RECT 106.53 12.19 106.77 13.06 ;
      RECT 106.95 14.52 107.11 16.86 ;
      RECT 106.82 13.22 106.98 14.84 ;
      RECT 106.55 41.08 106.71 45.17 ;
      RECT 106.55 41.08 106.87 41.24 ;
      RECT 105.73 17.6 105.89 23.81 ;
      RECT 105.25 22.38 106.37 22.54 ;
      RECT 105.73 58.24 105.89 64 ;
      RECT 105.25 59.51 106.37 59.67 ;
      RECT 106.15 27.37 106.31 31.49 ;
      RECT 105.31 27.37 105.47 31.49 ;
      RECT 105.31 27.37 106.31 27.53 ;
      RECT 105.73 24.64 105.89 27.53 ;
      RECT 105.73 54.16 105.89 57.42 ;
      RECT 105.31 54.16 106.31 54.88 ;
      RECT 106.15 50.8 106.31 54.88 ;
      RECT 105.31 50.8 105.47 54.88 ;
      RECT 103.57 55.09 104.83 55.25 ;
      RECT 104.67 49.77 104.83 55.25 ;
      RECT 104.67 49.77 105.55 49.93 ;
      RECT 105.39 32.48 105.55 49.93 ;
      RECT 104.73 45.9 105.55 46.06 ;
      RECT 104.73 36.23 105.55 36.39 ;
      RECT 104.67 32.48 105.55 32.64 ;
      RECT 104.67 27.04 104.83 32.64 ;
      RECT 103.57 27.04 104.83 27.2 ;
      RECT 103.47 26.46 105.49 26.62 ;
      RECT 105.33 25.35 105.49 26.62 ;
      RECT 105.25 22.91 105.41 25.51 ;
      RECT 105.25 56.46 105.41 59.14 ;
      RECT 105.33 55.49 105.49 56.62 ;
      RECT 103.47 55.49 105.49 55.65 ;
      RECT 102.82 71.82 103.1 72.56 ;
      RECT 102.82 71.87 105.37 72.42 ;
      RECT 103.49 71.86 105.37 72.42 ;
      RECT 104.93 25.79 105.17 26.07 ;
      RECT 104.93 21.94 105.09 26.07 ;
      RECT 104.93 21.94 105.21 22.18 ;
      RECT 104.99 15.28 105.15 22.18 ;
      RECT 104.03 15.28 104.19 20.88 ;
      RECT 103.07 15.28 103.23 20.88 ;
      RECT 103.07 17.14 105.15 17.3 ;
      RECT 104.99 59.87 105.15 66.77 ;
      RECT 104.03 61.17 104.19 66.77 ;
      RECT 103.07 61.17 103.23 66.77 ;
      RECT 103.07 64.75 105.15 64.91 ;
      RECT 104.93 59.87 105.21 60.11 ;
      RECT 104.93 56.02 105.09 60.11 ;
      RECT 104.93 56.02 105.17 56.3 ;
      RECT 103.07 35.91 105.15 36.07 ;
      RECT 104.99 32.85 105.15 36.07 ;
      RECT 104.03 27.43 104.19 36.07 ;
      RECT 103.07 32.85 103.23 36.07 ;
      RECT 103.13 27.43 104.19 27.59 ;
      RECT 103.13 23.41 103.29 27.59 ;
      RECT 103.13 26.14 104.29 26.3 ;
      RECT 104.13 25.01 104.29 26.3 ;
      RECT 103.13 25 103.33 26.3 ;
      RECT 104.13 21.38 104.29 23.81 ;
      RECT 103.17 21.38 103.33 23.55 ;
      RECT 103.17 21.38 104.29 21.54 ;
      RECT 103.17 60.51 104.29 60.67 ;
      RECT 104.13 58.24 104.29 60.67 ;
      RECT 103.17 58.5 103.33 60.67 ;
      RECT 103.13 55.81 103.29 58.64 ;
      RECT 104.13 55.81 104.29 57.09 ;
      RECT 103.11 55.81 103.33 57.09 ;
      RECT 103.11 55.81 104.29 55.97 ;
      RECT 103.11 54.64 103.27 57.09 ;
      RECT 103.11 54.64 104.19 54.8 ;
      RECT 104.03 46.22 104.19 54.8 ;
      RECT 104.99 46.22 105.15 49.44 ;
      RECT 103.07 46.22 103.23 49.44 ;
      RECT 103.07 46.22 105.15 46.38 ;
      RECT 104.43 12.8 105.09 13.06 ;
      RECT 104.85 12.19 105.09 13.06 ;
      RECT 104.91 41.08 105.07 45.17 ;
      RECT 104.75 41.08 105.07 41.24 ;
      RECT 104.61 21.06 104.77 26.28 ;
      RECT 103.65 24.37 103.81 25.98 ;
      RECT 103.45 24.37 104.77 24.53 ;
      RECT 103.45 23.67 103.61 24.53 ;
      RECT 103.45 23.67 103.81 23.83 ;
      RECT 103.65 21.7 103.81 23.83 ;
      RECT 102.95 21.06 104.83 21.22 ;
      RECT 102.95 60.83 104.83 60.99 ;
      RECT 104.61 55.81 104.77 60.99 ;
      RECT 103.65 58.22 103.81 60.35 ;
      RECT 103.45 58.22 103.81 58.38 ;
      RECT 103.45 57.25 103.61 58.38 ;
      RECT 103.45 57.25 104.77 57.41 ;
      RECT 103.65 56.13 103.81 57.41 ;
      RECT 104.51 14.52 104.67 16.86 ;
      RECT 104.64 13.22 104.8 14.84 ;
      RECT 104.51 32.85 104.67 35.75 ;
      RECT 104.35 31.09 104.51 33.01 ;
      RECT 104.35 49.44 104.51 51.3 ;
      RECT 104.51 46.54 104.67 49.6 ;
      RECT 104.43 38.57 104.59 45.17 ;
      RECT 104.13 38.57 104.59 38.73 ;
      RECT 104.13 36.23 104.29 38.73 ;
      RECT 103.77 36.23 104.45 36.39 ;
      RECT 103.65 45.9 104.45 46.06 ;
      RECT 103.65 44.89 103.81 46.06 ;
      RECT 103.63 38.57 103.79 45.17 ;
      RECT 104.03 10.09 104.19 14.2 ;
      RECT 103.13 12.9 104.19 13.06 ;
      RECT 103.13 12.19 103.29 13.06 ;
      RECT 103.55 14.52 103.71 16.86 ;
      RECT 103.42 13.22 103.58 14.84 ;
      RECT 103.55 31.09 103.71 35.75 ;
      RECT 103.45 32.25 103.71 32.53 ;
      RECT 103.51 49.75 103.71 51.3 ;
      RECT 103.55 46.54 103.71 51.3 ;
      RECT 103.11 49.6 103.27 51.7 ;
      RECT 102.67 49.6 103.27 49.76 ;
      RECT 102.67 32.06 102.83 49.76 ;
      RECT 102.67 45.9 103.49 46.06 ;
      RECT 102.67 36.23 103.49 36.39 ;
      RECT 102.67 32.06 103.27 32.22 ;
      RECT 103.11 30.54 103.27 32.22 ;
      RECT 103.15 41.08 103.31 45.17 ;
      RECT 103.15 41.08 103.47 41.24 ;
      RECT 102.33 31.49 102.49 32.02 ;
      RECT 101.87 31.49 102.95 31.65 ;
      RECT 102.79 27.38 102.95 31.65 ;
      RECT 101.87 27.38 102.03 31.65 ;
      RECT 101.87 27.38 102.95 27.54 ;
      RECT 102.33 26.91 102.49 27.54 ;
      RECT 101.87 51.06 102.95 55.29 ;
      RECT 102.33 50.27 102.49 55.29 ;
      RECT 102.69 49.92 102.85 50.9 ;
      RECT 101.97 49.92 102.13 50.9 ;
      RECT 101.97 49.92 102.85 50.08 ;
      RECT 102.33 45.65 102.49 50.08 ;
      RECT 101.55 49.6 101.71 51.7 ;
      RECT 101.55 49.6 102.15 49.76 ;
      RECT 101.99 32.06 102.15 49.76 ;
      RECT 101.33 45.9 102.15 46.06 ;
      RECT 101.33 36.23 102.15 36.39 ;
      RECT 101.55 32.06 102.15 32.22 ;
      RECT 101.55 30.54 101.71 32.22 ;
      RECT 99.42 71.82 99.7 72.56 ;
      RECT 99.42 71.87 101.97 72.42 ;
      RECT 100.09 71.86 101.97 72.42 ;
      RECT 99.42 85.42 99.7 86.16 ;
      RECT 99.42 85.47 101.97 86.02 ;
      RECT 100.09 85.46 101.97 86.02 ;
      RECT 99.42 99.02 99.7 99.76 ;
      RECT 99.42 99.07 101.97 99.62 ;
      RECT 100.09 99.06 101.97 99.62 ;
      RECT 99.42 112.62 99.7 113.36 ;
      RECT 99.42 112.67 101.97 113.22 ;
      RECT 100.09 112.66 101.97 113.22 ;
      RECT 99.42 126.22 99.7 126.96 ;
      RECT 99.42 126.27 101.97 126.82 ;
      RECT 100.09 126.26 101.97 126.82 ;
      RECT 99.42 139.82 99.7 140.56 ;
      RECT 99.42 139.87 101.97 140.42 ;
      RECT 100.09 139.86 101.97 140.42 ;
      RECT 99.42 153.42 99.7 154.16 ;
      RECT 99.42 153.47 101.97 154.02 ;
      RECT 100.09 153.46 101.97 154.02 ;
      RECT 99.42 167.02 99.7 167.76 ;
      RECT 99.42 167.07 101.97 167.62 ;
      RECT 100.09 167.06 101.97 167.62 ;
      RECT 99.42 180.62 99.7 181.36 ;
      RECT 99.42 180.67 101.97 181.22 ;
      RECT 100.09 180.66 101.97 181.22 ;
      RECT 99.42 194.22 99.7 194.96 ;
      RECT 99.42 194.27 101.97 194.82 ;
      RECT 100.09 194.26 101.97 194.82 ;
      RECT 99.42 207.82 99.7 208.56 ;
      RECT 99.42 207.87 101.97 208.42 ;
      RECT 100.09 207.86 101.97 208.42 ;
      RECT 99.42 221.42 99.7 222.16 ;
      RECT 99.42 221.47 101.97 222.02 ;
      RECT 100.09 221.46 101.97 222.02 ;
      RECT 99.42 235.02 99.7 235.76 ;
      RECT 99.42 235.07 101.97 235.62 ;
      RECT 100.09 235.06 101.97 235.62 ;
      RECT 99.42 248.62 99.7 249.36 ;
      RECT 99.42 248.67 101.97 249.22 ;
      RECT 100.09 248.66 101.97 249.22 ;
      RECT 99.42 262.22 99.7 262.96 ;
      RECT 99.42 262.27 101.97 262.82 ;
      RECT 100.09 262.26 101.97 262.82 ;
      RECT 99.42 275.82 99.7 276.56 ;
      RECT 99.42 275.87 101.97 276.42 ;
      RECT 100.09 275.86 101.97 276.42 ;
      RECT 99.42 289.42 99.7 290.16 ;
      RECT 99.42 289.47 101.97 290.02 ;
      RECT 100.09 289.46 101.97 290.02 ;
      RECT 99.42 303.02 99.7 303.76 ;
      RECT 99.42 303.07 101.97 303.62 ;
      RECT 100.09 303.06 101.97 303.62 ;
      RECT 99.42 316.62 99.7 317.36 ;
      RECT 99.42 316.67 101.97 317.22 ;
      RECT 100.09 316.66 101.97 317.22 ;
      RECT 99.42 330.22 99.7 330.96 ;
      RECT 99.42 330.27 101.97 330.82 ;
      RECT 100.09 330.26 101.97 330.82 ;
      RECT 99.42 343.82 99.7 344.56 ;
      RECT 99.42 343.87 101.97 344.42 ;
      RECT 100.09 343.86 101.97 344.42 ;
      RECT 99.42 357.42 99.7 358.16 ;
      RECT 99.42 357.47 101.97 358.02 ;
      RECT 100.09 357.46 101.97 358.02 ;
      RECT 99.42 371.02 99.7 371.76 ;
      RECT 99.42 371.07 101.97 371.62 ;
      RECT 100.09 371.06 101.97 371.62 ;
      RECT 99.42 384.62 99.7 385.36 ;
      RECT 99.42 384.67 101.97 385.22 ;
      RECT 100.09 384.66 101.97 385.22 ;
      RECT 99.42 398.22 99.7 398.96 ;
      RECT 99.42 398.27 101.97 398.82 ;
      RECT 100.09 398.26 101.97 398.82 ;
      RECT 99.42 411.82 99.7 412.56 ;
      RECT 99.42 411.87 101.97 412.42 ;
      RECT 100.09 411.86 101.97 412.42 ;
      RECT 99.42 425.42 99.7 426.16 ;
      RECT 99.42 425.47 101.97 426.02 ;
      RECT 100.09 425.46 101.97 426.02 ;
      RECT 99.42 439.02 99.7 439.76 ;
      RECT 99.42 439.07 101.97 439.62 ;
      RECT 100.09 439.06 101.97 439.62 ;
      RECT 99.42 452.62 99.7 453.36 ;
      RECT 99.42 452.67 101.97 453.22 ;
      RECT 100.09 452.66 101.97 453.22 ;
      RECT 99.42 466.22 99.7 466.96 ;
      RECT 99.42 466.27 101.97 466.82 ;
      RECT 100.09 466.26 101.97 466.82 ;
      RECT 99.42 479.82 99.7 480.56 ;
      RECT 99.42 479.87 101.97 480.42 ;
      RECT 100.09 479.86 101.97 480.42 ;
      RECT 99.42 493.42 99.7 494.16 ;
      RECT 99.42 493.47 101.97 494.02 ;
      RECT 100.09 493.46 101.97 494.02 ;
      RECT 100.05 21.06 100.21 26.28 ;
      RECT 101.01 24.37 101.17 25.98 ;
      RECT 100.05 24.37 101.37 24.53 ;
      RECT 101.21 23.67 101.37 24.53 ;
      RECT 101.01 23.67 101.37 23.83 ;
      RECT 101.01 21.7 101.17 23.83 ;
      RECT 99.99 21.06 101.87 21.22 ;
      RECT 99.99 60.83 101.87 60.99 ;
      RECT 100.05 55.81 100.21 60.99 ;
      RECT 101.01 58.22 101.17 60.35 ;
      RECT 101.01 58.22 101.37 58.38 ;
      RECT 101.21 57.25 101.37 58.38 ;
      RECT 100.05 57.25 101.37 57.41 ;
      RECT 101.01 56.13 101.17 57.41 ;
      RECT 99.65 25.79 99.89 26.07 ;
      RECT 99.73 21.94 99.89 26.07 ;
      RECT 99.61 21.94 99.89 22.18 ;
      RECT 99.67 15.28 99.83 22.18 ;
      RECT 101.59 15.28 101.75 20.88 ;
      RECT 100.63 15.28 100.79 20.88 ;
      RECT 99.67 17.14 101.75 17.3 ;
      RECT 99.67 35.91 101.75 36.07 ;
      RECT 101.59 32.85 101.75 36.07 ;
      RECT 100.63 27.43 100.79 36.07 ;
      RECT 99.67 32.85 99.83 36.07 ;
      RECT 100.63 27.43 101.69 27.59 ;
      RECT 101.53 23.41 101.69 27.59 ;
      RECT 100.53 26.14 101.69 26.3 ;
      RECT 101.49 25 101.69 26.3 ;
      RECT 100.53 25.01 100.69 26.3 ;
      RECT 100.53 21.38 100.69 23.81 ;
      RECT 101.49 21.38 101.65 23.55 ;
      RECT 100.53 21.38 101.65 21.54 ;
      RECT 100.53 60.51 101.65 60.67 ;
      RECT 101.49 58.5 101.65 60.67 ;
      RECT 101.53 55.81 101.65 60.67 ;
      RECT 100.53 58.24 100.69 60.67 ;
      RECT 101.55 54.64 101.69 58.64 ;
      RECT 101.49 55.81 101.71 57.09 ;
      RECT 101.55 54.64 101.71 57.09 ;
      RECT 100.53 55.81 100.69 57.09 ;
      RECT 100.53 55.81 101.71 55.97 ;
      RECT 100.63 54.64 101.71 54.8 ;
      RECT 100.63 46.22 100.79 54.8 ;
      RECT 101.59 46.22 101.75 49.44 ;
      RECT 99.67 46.22 99.83 49.44 ;
      RECT 99.67 46.22 101.75 46.38 ;
      RECT 101.59 61.17 101.75 66.77 ;
      RECT 100.63 61.17 100.79 66.77 ;
      RECT 99.67 59.87 99.83 66.77 ;
      RECT 99.67 64.75 101.75 64.91 ;
      RECT 99.61 59.87 99.89 60.11 ;
      RECT 99.73 56.02 99.89 60.11 ;
      RECT 99.65 56.02 99.89 56.3 ;
      RECT 100.63 10.09 100.79 14.2 ;
      RECT 100.63 12.9 101.69 13.06 ;
      RECT 101.53 12.19 101.69 13.06 ;
      RECT 101.51 41.08 101.67 45.17 ;
      RECT 101.35 41.08 101.67 41.24 ;
      RECT 101.11 14.52 101.27 16.86 ;
      RECT 101.24 13.22 101.4 14.84 ;
      RECT 101.11 31.09 101.27 35.75 ;
      RECT 101.11 32.25 101.37 32.53 ;
      RECT 99.33 26.46 101.35 26.62 ;
      RECT 99.33 25.35 99.49 26.62 ;
      RECT 99.41 22.91 99.57 25.51 ;
      RECT 99.41 56.46 99.57 59.14 ;
      RECT 99.33 55.49 99.49 56.62 ;
      RECT 99.33 55.49 101.35 55.65 ;
      RECT 101.11 49.75 101.31 51.3 ;
      RECT 101.11 46.54 101.27 51.3 ;
      RECT 99.99 55.09 101.25 55.25 ;
      RECT 99.99 49.77 100.15 55.25 ;
      RECT 99.27 49.77 100.15 49.93 ;
      RECT 99.27 32.48 99.43 49.93 ;
      RECT 99.27 45.9 100.09 46.06 ;
      RECT 99.27 36.23 100.09 36.39 ;
      RECT 99.27 32.48 100.15 32.64 ;
      RECT 99.99 27.04 100.15 32.64 ;
      RECT 99.99 27.04 101.25 27.2 ;
      RECT 100.37 45.9 101.17 46.06 ;
      RECT 101.01 44.89 101.17 46.06 ;
      RECT 101.03 38.57 101.19 45.17 ;
      RECT 100.23 38.57 100.39 45.17 ;
      RECT 100.23 38.57 100.69 38.73 ;
      RECT 100.53 36.23 100.69 38.73 ;
      RECT 100.37 36.23 101.05 36.39 ;
      RECT 100.15 32.85 100.31 35.75 ;
      RECT 100.31 31.09 100.47 33.01 ;
      RECT 100.31 49.44 100.47 51.3 ;
      RECT 100.15 46.54 100.31 49.6 ;
      RECT 99.73 12.8 100.39 13.06 ;
      RECT 99.73 12.19 99.97 13.06 ;
      RECT 100.15 14.52 100.31 16.86 ;
      RECT 100.02 13.22 100.18 14.84 ;
      RECT 99.75 41.08 99.91 45.17 ;
      RECT 99.75 41.08 100.07 41.24 ;
      RECT 98.93 17.6 99.09 23.81 ;
      RECT 98.45 22.38 99.57 22.54 ;
      RECT 98.93 58.24 99.09 64 ;
      RECT 98.45 59.51 99.57 59.67 ;
      RECT 99.35 27.37 99.51 31.49 ;
      RECT 98.51 27.37 98.67 31.49 ;
      RECT 98.51 27.37 99.51 27.53 ;
      RECT 98.93 24.64 99.09 27.53 ;
      RECT 98.93 54.16 99.09 57.42 ;
      RECT 98.51 54.16 99.51 54.88 ;
      RECT 99.35 50.8 99.51 54.88 ;
      RECT 98.51 50.8 98.67 54.88 ;
      RECT 96.77 55.09 98.03 55.25 ;
      RECT 97.87 49.77 98.03 55.25 ;
      RECT 97.87 49.77 98.75 49.93 ;
      RECT 98.59 32.48 98.75 49.93 ;
      RECT 97.93 45.9 98.75 46.06 ;
      RECT 97.93 36.23 98.75 36.39 ;
      RECT 97.87 32.48 98.75 32.64 ;
      RECT 97.87 27.04 98.03 32.64 ;
      RECT 96.77 27.04 98.03 27.2 ;
      RECT 96.67 26.46 98.69 26.62 ;
      RECT 98.53 25.35 98.69 26.62 ;
      RECT 98.45 22.91 98.61 25.51 ;
      RECT 98.45 56.46 98.61 59.14 ;
      RECT 98.53 55.49 98.69 56.62 ;
      RECT 96.67 55.49 98.69 55.65 ;
      RECT 98.04 9.18 98.2 14.23 ;
      RECT 96.51 9.18 96.67 14.23 ;
      RECT 96.51 11.85 98.2 12.01 ;
      RECT 96.51 9.18 98.2 9.34 ;
      RECT 96.98 7.64 97.66 9.34 ;
      RECT 96.25 7.64 98.53 8.28 ;
      RECT 98.13 25.79 98.37 26.07 ;
      RECT 98.13 21.94 98.29 26.07 ;
      RECT 98.13 21.94 98.41 22.18 ;
      RECT 98.19 15.28 98.35 22.18 ;
      RECT 97.23 15.28 97.39 20.88 ;
      RECT 96.27 15.28 96.43 20.88 ;
      RECT 96.27 17.14 98.35 17.3 ;
      RECT 98.19 59.87 98.35 66.77 ;
      RECT 97.23 61.17 97.39 66.77 ;
      RECT 96.27 61.17 96.43 66.77 ;
      RECT 96.27 64.75 98.35 64.91 ;
      RECT 98.13 59.87 98.41 60.11 ;
      RECT 98.13 56.02 98.29 60.11 ;
      RECT 98.13 56.02 98.37 56.3 ;
      RECT 96.02 71.82 96.3 72.56 ;
      RECT 96.03 69.79 96.19 72.56 ;
      RECT 96.03 71.33 98.4 71.49 ;
      RECT 96.03 69.79 98.4 69.95 ;
      RECT 96.02 85.42 96.3 86.16 ;
      RECT 96.03 83.39 96.19 86.16 ;
      RECT 96.03 84.93 98.4 85.09 ;
      RECT 96.03 83.39 98.4 83.55 ;
      RECT 96.02 99.02 96.3 99.76 ;
      RECT 96.03 96.99 96.19 99.76 ;
      RECT 96.03 98.53 98.4 98.69 ;
      RECT 96.03 96.99 98.4 97.15 ;
      RECT 96.02 112.62 96.3 113.36 ;
      RECT 96.03 110.59 96.19 113.36 ;
      RECT 96.03 112.13 98.4 112.29 ;
      RECT 96.03 110.59 98.4 110.75 ;
      RECT 96.02 126.22 96.3 126.96 ;
      RECT 96.03 124.19 96.19 126.96 ;
      RECT 96.03 125.73 98.4 125.89 ;
      RECT 96.03 124.19 98.4 124.35 ;
      RECT 96.02 139.82 96.3 140.56 ;
      RECT 96.03 137.79 96.19 140.56 ;
      RECT 96.03 139.33 98.4 139.49 ;
      RECT 96.03 137.79 98.4 137.95 ;
      RECT 96.02 153.42 96.3 154.16 ;
      RECT 96.03 151.39 96.19 154.16 ;
      RECT 96.03 152.93 98.4 153.09 ;
      RECT 96.03 151.39 98.4 151.55 ;
      RECT 96.02 167.02 96.3 167.76 ;
      RECT 96.03 164.99 96.19 167.76 ;
      RECT 96.03 166.53 98.4 166.69 ;
      RECT 96.03 164.99 98.4 165.15 ;
      RECT 96.02 180.62 96.3 181.36 ;
      RECT 96.03 178.59 96.19 181.36 ;
      RECT 96.03 180.13 98.4 180.29 ;
      RECT 96.03 178.59 98.4 178.75 ;
      RECT 96.02 194.22 96.3 194.96 ;
      RECT 96.03 192.19 96.19 194.96 ;
      RECT 96.03 193.73 98.4 193.89 ;
      RECT 96.03 192.19 98.4 192.35 ;
      RECT 96.02 207.82 96.3 208.56 ;
      RECT 96.03 205.79 96.19 208.56 ;
      RECT 96.03 207.33 98.4 207.49 ;
      RECT 96.03 205.79 98.4 205.95 ;
      RECT 96.02 221.42 96.3 222.16 ;
      RECT 96.03 219.39 96.19 222.16 ;
      RECT 96.03 220.93 98.4 221.09 ;
      RECT 96.03 219.39 98.4 219.55 ;
      RECT 96.02 235.02 96.3 235.76 ;
      RECT 96.03 232.99 96.19 235.76 ;
      RECT 96.03 234.53 98.4 234.69 ;
      RECT 96.03 232.99 98.4 233.15 ;
      RECT 96.02 248.62 96.3 249.36 ;
      RECT 96.03 246.59 96.19 249.36 ;
      RECT 96.03 248.13 98.4 248.29 ;
      RECT 96.03 246.59 98.4 246.75 ;
      RECT 96.02 262.22 96.3 262.96 ;
      RECT 96.03 260.19 96.19 262.96 ;
      RECT 96.03 261.73 98.4 261.89 ;
      RECT 96.03 260.19 98.4 260.35 ;
      RECT 96.02 275.82 96.3 276.56 ;
      RECT 96.03 273.79 96.19 276.56 ;
      RECT 96.03 275.33 98.4 275.49 ;
      RECT 96.03 273.79 98.4 273.95 ;
      RECT 96.02 289.42 96.3 290.16 ;
      RECT 96.03 287.39 96.19 290.16 ;
      RECT 96.03 288.93 98.4 289.09 ;
      RECT 96.03 287.39 98.4 287.55 ;
      RECT 96.02 303.02 96.3 303.76 ;
      RECT 96.03 300.99 96.19 303.76 ;
      RECT 96.03 302.53 98.4 302.69 ;
      RECT 96.03 300.99 98.4 301.15 ;
      RECT 96.02 316.62 96.3 317.36 ;
      RECT 96.03 314.59 96.19 317.36 ;
      RECT 96.03 316.13 98.4 316.29 ;
      RECT 96.03 314.59 98.4 314.75 ;
      RECT 96.02 330.22 96.3 330.96 ;
      RECT 96.03 328.19 96.19 330.96 ;
      RECT 96.03 329.73 98.4 329.89 ;
      RECT 96.03 328.19 98.4 328.35 ;
      RECT 96.02 343.82 96.3 344.56 ;
      RECT 96.03 341.79 96.19 344.56 ;
      RECT 96.03 343.33 98.4 343.49 ;
      RECT 96.03 341.79 98.4 341.95 ;
      RECT 96.02 357.42 96.3 358.16 ;
      RECT 96.03 355.39 96.19 358.16 ;
      RECT 96.03 356.93 98.4 357.09 ;
      RECT 96.03 355.39 98.4 355.55 ;
      RECT 96.02 371.02 96.3 371.76 ;
      RECT 96.03 368.99 96.19 371.76 ;
      RECT 96.03 370.53 98.4 370.69 ;
      RECT 96.03 368.99 98.4 369.15 ;
      RECT 96.02 384.62 96.3 385.36 ;
      RECT 96.03 382.59 96.19 385.36 ;
      RECT 96.03 384.13 98.4 384.29 ;
      RECT 96.03 382.59 98.4 382.75 ;
      RECT 96.02 398.22 96.3 398.96 ;
      RECT 96.03 396.19 96.19 398.96 ;
      RECT 96.03 397.73 98.4 397.89 ;
      RECT 96.03 396.19 98.4 396.35 ;
      RECT 96.02 411.82 96.3 412.56 ;
      RECT 96.03 409.79 96.19 412.56 ;
      RECT 96.03 411.33 98.4 411.49 ;
      RECT 96.03 409.79 98.4 409.95 ;
      RECT 96.02 425.42 96.3 426.16 ;
      RECT 96.03 423.39 96.19 426.16 ;
      RECT 96.03 424.93 98.4 425.09 ;
      RECT 96.03 423.39 98.4 423.55 ;
      RECT 96.02 439.02 96.3 439.76 ;
      RECT 96.03 436.99 96.19 439.76 ;
      RECT 96.03 438.53 98.4 438.69 ;
      RECT 96.03 436.99 98.4 437.15 ;
      RECT 96.02 452.62 96.3 453.36 ;
      RECT 96.03 450.59 96.19 453.36 ;
      RECT 96.03 452.13 98.4 452.29 ;
      RECT 96.03 450.59 98.4 450.75 ;
      RECT 96.02 466.22 96.3 466.96 ;
      RECT 96.03 464.19 96.19 466.96 ;
      RECT 96.03 465.73 98.4 465.89 ;
      RECT 96.03 464.19 98.4 464.35 ;
      RECT 96.02 479.82 96.3 480.56 ;
      RECT 96.03 477.79 96.19 480.56 ;
      RECT 96.03 479.33 98.4 479.49 ;
      RECT 96.03 477.79 98.4 477.95 ;
      RECT 96.02 493.42 96.3 494.16 ;
      RECT 96.03 491.39 96.19 494.16 ;
      RECT 96.03 492.93 98.4 493.09 ;
      RECT 96.03 491.39 98.4 491.55 ;
      RECT 96.27 35.91 98.35 36.07 ;
      RECT 98.19 32.85 98.35 36.07 ;
      RECT 97.23 27.43 97.39 36.07 ;
      RECT 96.27 32.85 96.43 36.07 ;
      RECT 96.33 27.43 97.39 27.59 ;
      RECT 96.33 23.41 96.49 27.59 ;
      RECT 96.33 26.14 97.49 26.3 ;
      RECT 97.33 25.01 97.49 26.3 ;
      RECT 96.33 25 96.53 26.3 ;
      RECT 97.33 21.38 97.49 23.81 ;
      RECT 96.37 21.38 96.53 23.55 ;
      RECT 96.37 21.38 97.49 21.54 ;
      RECT 96.37 60.51 97.49 60.67 ;
      RECT 97.33 58.24 97.49 60.67 ;
      RECT 96.37 58.5 96.53 60.67 ;
      RECT 96.33 55.81 96.49 58.64 ;
      RECT 97.33 55.81 97.49 57.09 ;
      RECT 96.31 55.81 96.53 57.09 ;
      RECT 96.31 55.81 97.49 55.97 ;
      RECT 96.31 54.64 96.47 57.09 ;
      RECT 96.31 54.64 97.39 54.8 ;
      RECT 97.23 46.22 97.39 54.8 ;
      RECT 98.19 46.22 98.35 49.44 ;
      RECT 96.27 46.22 96.43 49.44 ;
      RECT 96.27 46.22 98.35 46.38 ;
      RECT 98.11 41.08 98.27 45.17 ;
      RECT 97.95 41.08 98.27 41.24 ;
      RECT 97.81 21.06 97.97 26.28 ;
      RECT 96.85 24.37 97.01 25.98 ;
      RECT 96.65 24.37 97.97 24.53 ;
      RECT 96.65 23.67 96.81 24.53 ;
      RECT 96.65 23.67 97.01 23.83 ;
      RECT 96.85 21.7 97.01 23.83 ;
      RECT 96.15 21.06 98.03 21.22 ;
      RECT 96.15 60.83 98.03 60.99 ;
      RECT 97.81 55.81 97.97 60.99 ;
      RECT 96.85 58.22 97.01 60.35 ;
      RECT 96.65 58.22 97.01 58.38 ;
      RECT 96.65 57.25 96.81 58.38 ;
      RECT 96.65 57.25 97.97 57.41 ;
      RECT 96.85 56.13 97.01 57.41 ;
      RECT 97.71 32.85 97.87 35.75 ;
      RECT 97.55 31.09 97.71 33.01 ;
      RECT 97.55 49.44 97.71 51.3 ;
      RECT 97.71 46.54 97.87 49.6 ;
      RECT 97.63 38.57 97.79 45.17 ;
      RECT 97.33 38.57 97.79 38.73 ;
      RECT 97.33 36.23 97.49 38.73 ;
      RECT 96.97 36.23 97.65 36.39 ;
      RECT 96.85 45.9 97.65 46.06 ;
      RECT 96.85 44.89 97.01 46.06 ;
      RECT 96.83 38.57 96.99 45.17 ;
      RECT 96.75 31.09 96.91 35.75 ;
      RECT 96.65 32.25 96.91 32.53 ;
      RECT 96.71 49.75 96.91 51.3 ;
      RECT 96.75 46.54 96.91 51.3 ;
      RECT 96.31 49.6 96.47 51.7 ;
      RECT 95.87 49.6 96.47 49.76 ;
      RECT 95.87 32.06 96.03 49.76 ;
      RECT 95.87 45.9 96.69 46.06 ;
      RECT 95.87 36.23 96.69 36.39 ;
      RECT 95.87 32.06 96.47 32.22 ;
      RECT 96.31 30.54 96.47 32.22 ;
      RECT 96.35 41.08 96.51 45.17 ;
      RECT 96.35 41.08 96.67 41.24 ;
      RECT 95.53 31.49 95.69 32.02 ;
      RECT 95.07 31.49 96.15 31.65 ;
      RECT 95.99 27.38 96.15 31.65 ;
      RECT 95.07 27.38 95.23 31.65 ;
      RECT 95.07 27.38 96.15 27.54 ;
      RECT 95.53 26.91 95.69 27.54 ;
      RECT 95.07 51.06 96.15 55.29 ;
      RECT 95.53 50.27 95.69 55.29 ;
      RECT 95.89 49.92 96.05 50.9 ;
      RECT 95.17 49.92 95.33 50.9 ;
      RECT 95.17 49.92 96.05 50.08 ;
      RECT 95.53 45.65 95.69 50.08 ;
      RECT 94.27 12.34 94.55 12.62 ;
      RECT 93.35 12.34 93.63 12.62 ;
      RECT 90.79 12.34 91.07 12.62 ;
      RECT 89.87 12.34 90.15 12.62 ;
      RECT 94.39 11.75 94.55 12.62 ;
      RECT 93.35 11.75 93.51 12.62 ;
      RECT 90.91 11.75 91.07 12.62 ;
      RECT 89.87 11.75 90.03 12.62 ;
      RECT 95.53 8.38 95.69 12.03 ;
      RECT 94.43 9.02 94.59 12.03 ;
      RECT 93.23 9.02 93.39 12.03 ;
      RECT 92.13 8.38 92.29 12.03 ;
      RECT 91.03 9.02 91.19 12.03 ;
      RECT 89.83 9.02 89.99 12.03 ;
      RECT 88.73 8.38 88.89 12.03 ;
      RECT 88.73 9.02 95.69 9.3 ;
      RECT 94.85 8.38 95.09 9.3 ;
      RECT 94.17 8.38 94.41 9.3 ;
      RECT 93.42 8.38 93.66 9.3 ;
      RECT 92.73 8.38 92.97 9.3 ;
      RECT 91.45 8.38 91.69 9.3 ;
      RECT 90.76 8.38 91 9.3 ;
      RECT 90.01 8.38 90.25 9.3 ;
      RECT 89.33 8.38 89.57 9.3 ;
      RECT 94.75 49.6 94.91 51.7 ;
      RECT 94.75 49.6 95.35 49.76 ;
      RECT 95.19 32.06 95.35 49.76 ;
      RECT 94.53 45.9 95.35 46.06 ;
      RECT 94.53 36.23 95.35 36.39 ;
      RECT 94.75 32.06 95.35 32.22 ;
      RECT 94.75 30.54 94.91 32.22 ;
      RECT 93.25 21.06 93.41 26.28 ;
      RECT 94.21 24.37 94.37 25.98 ;
      RECT 93.25 24.37 94.57 24.53 ;
      RECT 94.41 23.67 94.57 24.53 ;
      RECT 94.21 23.67 94.57 23.83 ;
      RECT 94.21 21.7 94.37 23.83 ;
      RECT 93.19 21.06 95.07 21.22 ;
      RECT 93.19 60.83 95.07 60.99 ;
      RECT 93.25 55.81 93.41 60.99 ;
      RECT 94.21 58.22 94.37 60.35 ;
      RECT 94.21 58.22 94.57 58.38 ;
      RECT 94.41 57.25 94.57 58.38 ;
      RECT 93.25 57.25 94.57 57.41 ;
      RECT 94.21 56.13 94.37 57.41 ;
      RECT 92.85 25.79 93.09 26.07 ;
      RECT 92.93 21.94 93.09 26.07 ;
      RECT 92.81 21.94 93.09 22.18 ;
      RECT 92.87 15.28 93.03 22.18 ;
      RECT 94.79 15.28 94.95 20.88 ;
      RECT 93.83 15.28 93.99 20.88 ;
      RECT 92.87 17.14 94.95 17.3 ;
      RECT 92.87 35.91 94.95 36.07 ;
      RECT 94.79 32.85 94.95 36.07 ;
      RECT 93.83 27.43 93.99 36.07 ;
      RECT 92.87 32.85 93.03 36.07 ;
      RECT 93.83 27.43 94.89 27.59 ;
      RECT 94.73 23.41 94.89 27.59 ;
      RECT 93.73 26.14 94.89 26.3 ;
      RECT 94.69 25 94.89 26.3 ;
      RECT 93.73 25.01 93.89 26.3 ;
      RECT 93.73 21.38 93.89 23.81 ;
      RECT 94.69 21.38 94.85 23.55 ;
      RECT 93.73 21.38 94.85 21.54 ;
      RECT 93.73 60.51 94.85 60.67 ;
      RECT 94.69 58.5 94.85 60.67 ;
      RECT 94.73 55.81 94.85 60.67 ;
      RECT 93.73 58.24 93.89 60.67 ;
      RECT 94.75 54.64 94.89 58.64 ;
      RECT 94.69 55.81 94.91 57.09 ;
      RECT 94.75 54.64 94.91 57.09 ;
      RECT 93.73 55.81 93.89 57.09 ;
      RECT 93.73 55.81 94.91 55.97 ;
      RECT 93.83 54.64 94.91 54.8 ;
      RECT 93.83 46.22 93.99 54.8 ;
      RECT 94.79 46.22 94.95 49.44 ;
      RECT 92.87 46.22 93.03 49.44 ;
      RECT 92.87 46.22 94.95 46.38 ;
      RECT 94.79 61.17 94.95 66.77 ;
      RECT 93.83 61.17 93.99 66.77 ;
      RECT 92.87 59.87 93.03 66.77 ;
      RECT 92.87 64.75 94.95 64.91 ;
      RECT 92.81 59.87 93.09 60.11 ;
      RECT 92.93 56.02 93.09 60.11 ;
      RECT 92.85 56.02 93.09 56.3 ;
      RECT 93.83 10.09 93.99 14.2 ;
      RECT 93.83 12.9 94.89 13.06 ;
      RECT 94.73 12.19 94.89 13.06 ;
      RECT 94.71 41.08 94.87 45.17 ;
      RECT 94.55 41.08 94.87 41.24 ;
      RECT 94.31 14.52 94.47 16.86 ;
      RECT 94.44 13.22 94.6 14.84 ;
      RECT 94.31 31.09 94.47 35.75 ;
      RECT 94.31 32.25 94.57 32.53 ;
      RECT 92.53 26.46 94.55 26.62 ;
      RECT 92.53 25.35 92.69 26.62 ;
      RECT 92.61 22.91 92.77 25.51 ;
      RECT 92.61 56.46 92.77 59.14 ;
      RECT 92.53 55.49 92.69 56.62 ;
      RECT 92.53 55.49 94.55 55.65 ;
      RECT 94.31 49.75 94.51 51.3 ;
      RECT 94.31 46.54 94.47 51.3 ;
      RECT 93.19 55.09 94.45 55.25 ;
      RECT 93.19 49.77 93.35 55.25 ;
      RECT 92.47 49.77 93.35 49.93 ;
      RECT 92.47 32.48 92.63 49.93 ;
      RECT 92.47 45.9 93.29 46.06 ;
      RECT 92.47 36.23 93.29 36.39 ;
      RECT 92.47 32.48 93.35 32.64 ;
      RECT 93.19 27.04 93.35 32.64 ;
      RECT 93.19 27.04 94.45 27.2 ;
      RECT 93.57 45.9 94.37 46.06 ;
      RECT 94.21 44.89 94.37 46.06 ;
      RECT 94.23 38.57 94.39 45.17 ;
      RECT 93.43 38.57 93.59 45.17 ;
      RECT 93.43 38.57 93.89 38.73 ;
      RECT 93.73 36.23 93.89 38.73 ;
      RECT 93.57 36.23 94.25 36.39 ;
      RECT 93.35 32.85 93.51 35.75 ;
      RECT 93.51 31.09 93.67 33.01 ;
      RECT 93.51 49.44 93.67 51.3 ;
      RECT 93.35 46.54 93.51 49.6 ;
      RECT 92.93 12.8 93.59 13.06 ;
      RECT 92.93 12.19 93.17 13.06 ;
      RECT 93.35 14.52 93.51 16.86 ;
      RECT 93.22 13.22 93.38 14.84 ;
      RECT 92.95 41.08 93.11 45.17 ;
      RECT 92.95 41.08 93.27 41.24 ;
      RECT 92.13 17.6 92.29 23.81 ;
      RECT 91.65 22.38 92.77 22.54 ;
      RECT 92.13 58.24 92.29 64 ;
      RECT 91.65 59.51 92.77 59.67 ;
      RECT 92.55 27.37 92.71 31.49 ;
      RECT 91.71 27.37 91.87 31.49 ;
      RECT 91.71 27.37 92.71 27.53 ;
      RECT 92.13 24.64 92.29 27.53 ;
      RECT 92.13 54.16 92.29 57.42 ;
      RECT 91.71 54.16 92.71 54.88 ;
      RECT 92.55 50.8 92.71 54.88 ;
      RECT 91.71 50.8 91.87 54.88 ;
      RECT 89.97 55.09 91.23 55.25 ;
      RECT 91.07 49.77 91.23 55.25 ;
      RECT 91.07 49.77 91.95 49.93 ;
      RECT 91.79 32.48 91.95 49.93 ;
      RECT 91.13 45.9 91.95 46.06 ;
      RECT 91.13 36.23 91.95 36.39 ;
      RECT 91.07 32.48 91.95 32.64 ;
      RECT 91.07 27.04 91.23 32.64 ;
      RECT 89.97 27.04 91.23 27.2 ;
      RECT 89.87 26.46 91.89 26.62 ;
      RECT 91.73 25.35 91.89 26.62 ;
      RECT 91.65 22.91 91.81 25.51 ;
      RECT 91.65 56.46 91.81 59.14 ;
      RECT 91.73 55.49 91.89 56.62 ;
      RECT 89.87 55.49 91.89 55.65 ;
      RECT 91.33 25.79 91.57 26.07 ;
      RECT 91.33 21.94 91.49 26.07 ;
      RECT 91.33 21.94 91.61 22.18 ;
      RECT 91.39 15.28 91.55 22.18 ;
      RECT 90.43 15.28 90.59 20.88 ;
      RECT 89.47 15.28 89.63 20.88 ;
      RECT 89.47 17.14 91.55 17.3 ;
      RECT 91.39 59.87 91.55 66.77 ;
      RECT 90.43 61.17 90.59 66.77 ;
      RECT 89.47 61.17 89.63 66.77 ;
      RECT 89.47 64.75 91.55 64.91 ;
      RECT 91.33 59.87 91.61 60.11 ;
      RECT 91.33 56.02 91.49 60.11 ;
      RECT 91.33 56.02 91.57 56.3 ;
      RECT 89.47 35.91 91.55 36.07 ;
      RECT 91.39 32.85 91.55 36.07 ;
      RECT 90.43 27.43 90.59 36.07 ;
      RECT 89.47 32.85 89.63 36.07 ;
      RECT 89.53 27.43 90.59 27.59 ;
      RECT 89.53 23.41 89.69 27.59 ;
      RECT 89.53 26.14 90.69 26.3 ;
      RECT 90.53 25.01 90.69 26.3 ;
      RECT 89.53 25 89.73 26.3 ;
      RECT 90.53 21.38 90.69 23.81 ;
      RECT 89.57 21.38 89.73 23.55 ;
      RECT 89.57 21.38 90.69 21.54 ;
      RECT 89.57 60.51 90.69 60.67 ;
      RECT 90.53 58.24 90.69 60.67 ;
      RECT 89.57 58.5 89.73 60.67 ;
      RECT 89.53 55.81 89.69 58.64 ;
      RECT 90.53 55.81 90.69 57.09 ;
      RECT 89.51 55.81 89.73 57.09 ;
      RECT 89.51 55.81 90.69 55.97 ;
      RECT 89.51 54.64 89.67 57.09 ;
      RECT 89.51 54.64 90.59 54.8 ;
      RECT 90.43 46.22 90.59 54.8 ;
      RECT 91.39 46.22 91.55 49.44 ;
      RECT 89.47 46.22 89.63 49.44 ;
      RECT 89.47 46.22 91.55 46.38 ;
      RECT 90.83 12.8 91.49 13.06 ;
      RECT 91.25 12.19 91.49 13.06 ;
      RECT 91.31 41.08 91.47 45.17 ;
      RECT 91.15 41.08 91.47 41.24 ;
      RECT 91.01 21.06 91.17 26.28 ;
      RECT 90.05 24.37 90.21 25.98 ;
      RECT 89.85 24.37 91.17 24.53 ;
      RECT 89.85 23.67 90.01 24.53 ;
      RECT 89.85 23.67 90.21 23.83 ;
      RECT 90.05 21.7 90.21 23.83 ;
      RECT 89.35 21.06 91.23 21.22 ;
      RECT 89.35 60.83 91.23 60.99 ;
      RECT 91.01 55.81 91.17 60.99 ;
      RECT 90.05 58.22 90.21 60.35 ;
      RECT 89.85 58.22 90.21 58.38 ;
      RECT 89.85 57.25 90.01 58.38 ;
      RECT 89.85 57.25 91.17 57.41 ;
      RECT 90.05 56.13 90.21 57.41 ;
      RECT 90.91 14.52 91.07 16.86 ;
      RECT 91.04 13.22 91.2 14.84 ;
      RECT 90.91 32.85 91.07 35.75 ;
      RECT 90.75 31.09 90.91 33.01 ;
      RECT 90.75 49.44 90.91 51.3 ;
      RECT 90.91 46.54 91.07 49.6 ;
      RECT 90.83 38.57 90.99 45.17 ;
      RECT 90.53 38.57 90.99 38.73 ;
      RECT 90.53 36.23 90.69 38.73 ;
      RECT 90.17 36.23 90.85 36.39 ;
      RECT 90.05 45.9 90.85 46.06 ;
      RECT 90.05 44.89 90.21 46.06 ;
      RECT 90.03 38.57 90.19 45.17 ;
      RECT 90.43 10.09 90.59 14.2 ;
      RECT 89.53 12.9 90.59 13.06 ;
      RECT 89.53 12.19 89.69 13.06 ;
      RECT 89.95 14.52 90.11 16.86 ;
      RECT 89.82 13.22 89.98 14.84 ;
      RECT 89.95 31.09 90.11 35.75 ;
      RECT 89.85 32.25 90.11 32.53 ;
      RECT 89.91 49.75 90.11 51.3 ;
      RECT 89.95 46.54 90.11 51.3 ;
      RECT 89.51 49.6 89.67 51.7 ;
      RECT 89.07 49.6 89.67 49.76 ;
      RECT 89.07 32.06 89.23 49.76 ;
      RECT 89.07 45.9 89.89 46.06 ;
      RECT 89.07 36.23 89.89 36.39 ;
      RECT 89.07 32.06 89.67 32.22 ;
      RECT 89.51 30.54 89.67 32.22 ;
      RECT 89.55 41.08 89.71 45.17 ;
      RECT 89.55 41.08 89.87 41.24 ;
      RECT 88.73 31.49 88.89 32.02 ;
      RECT 88.73 31.49 89.35 31.65 ;
      RECT 89.19 27.38 89.35 31.65 ;
      RECT 88.73 27.38 89.35 27.54 ;
      RECT 88.73 26.91 88.89 27.54 ;
      RECT 88.73 51.06 89.35 55.29 ;
      RECT 88.73 50.27 88.89 55.29 ;
      RECT 89.09 49.92 89.25 50.9 ;
      RECT 88.73 49.92 89.25 50.08 ;
      RECT 88.73 45.65 88.89 50.08 ;
      RECT 86.33 46.75 86.49 47.43 ;
      RECT 86.01 46.75 86.49 46.91 ;
      RECT 86.01 44.23 86.17 46.91 ;
      RECT 8.33 68.47 86.49 68.63 ;
      RECT 86.33 56.96 86.49 68.63 ;
      RECT 83.93 56.96 84.09 68.63 ;
      RECT 81.53 56.96 81.69 68.63 ;
      RECT 79.13 56.96 79.29 68.63 ;
      RECT 76.73 56.96 76.89 68.63 ;
      RECT 74.33 56.96 74.49 68.63 ;
      RECT 71.93 56.96 72.09 68.63 ;
      RECT 69.53 56.96 69.69 68.63 ;
      RECT 67.13 56.96 67.29 68.63 ;
      RECT 64.73 56.96 64.89 68.63 ;
      RECT 62.33 56.96 62.49 68.63 ;
      RECT 59.93 56.96 60.09 68.63 ;
      RECT 57.53 56.96 57.69 68.63 ;
      RECT 55.13 56.96 55.29 68.63 ;
      RECT 52.73 56.96 52.89 68.63 ;
      RECT 50.33 56.96 50.49 68.63 ;
      RECT 47.93 56.96 48.09 68.63 ;
      RECT 46.73 56.96 46.89 68.63 ;
      RECT 44.33 56.96 44.49 68.63 ;
      RECT 41.93 56.96 42.09 68.63 ;
      RECT 39.53 56.96 39.69 68.63 ;
      RECT 37.13 56.96 37.29 68.63 ;
      RECT 34.73 56.96 34.89 68.63 ;
      RECT 32.33 56.96 32.49 68.63 ;
      RECT 29.93 56.96 30.09 68.63 ;
      RECT 27.53 56.96 27.69 68.63 ;
      RECT 25.13 56.96 25.29 68.63 ;
      RECT 22.73 56.96 22.89 68.63 ;
      RECT 20.33 56.96 20.49 68.63 ;
      RECT 17.93 56.96 18.09 68.63 ;
      RECT 15.53 56.96 15.69 68.63 ;
      RECT 13.13 56.96 13.29 68.63 ;
      RECT 10.73 56.96 10.89 68.63 ;
      RECT 8.33 56.96 8.49 68.63 ;
      RECT 84.11 34.88 86.31 35.04 ;
      RECT 86.03 34.59 86.31 35.04 ;
      RECT 85.09 34.59 85.33 35.04 ;
      RECT 84.11 34.59 84.39 35.04 ;
      RECT 85.09 38.38 85.33 39.02 ;
      RECT 86.03 38.38 86.31 38.83 ;
      RECT 84.11 38.38 84.39 38.83 ;
      RECT 84.11 38.38 86.31 38.54 ;
      RECT 84.27 36.47 86.15 36.63 ;
      RECT 85.99 35.88 86.15 36.63 ;
      RECT 85.13 35.23 85.29 36.63 ;
      RECT 84.27 35.88 84.43 36.63 ;
      RECT 86.09 35.23 86.25 36.06 ;
      RECT 84.17 35.23 84.33 36.06 ;
      RECT 86.09 37.11 86.25 38.19 ;
      RECT 85.13 36.79 85.29 38.19 ;
      RECT 84.17 37.11 84.33 38.19 ;
      RECT 85.99 36.79 86.15 37.39 ;
      RECT 84.27 36.79 84.43 37.39 ;
      RECT 84.27 36.79 86.15 36.95 ;
      RECT 84.35 68.07 86.17 68.23 ;
      RECT 84.35 62.02 84.51 68.23 ;
      RECT 84.35 62.02 84.73 62.18 ;
      RECT 84.57 57.45 84.73 62.18 ;
      RECT 84.57 57.45 86.17 57.61 ;
      RECT 85.85 57.39 86.17 57.61 ;
      RECT 85.85 53.74 86.01 57.61 ;
      RECT 86.01 51.32 86.17 53.9 ;
      RECT 85.69 51.32 86.17 51.48 ;
      RECT 85.69 49.88 85.85 51.48 ;
      RECT 85.37 49.88 85.85 50.04 ;
      RECT 85.37 47.71 85.53 50.04 ;
      RECT 84.91 47.71 85.53 47.99 ;
      RECT 85.69 47.39 85.85 49.72 ;
      RECT 85.37 47.39 85.85 47.55 ;
      RECT 85.37 43.85 85.53 47.55 ;
      RECT 85.37 43.85 86.15 44.01 ;
      RECT 85.99 39.56 86.15 44.01 ;
      RECT 85.81 39.56 86.15 39.84 ;
      RECT 85.81 39.16 85.97 39.84 ;
      RECT 85.85 62.9 86.01 67.89 ;
      RECT 85.73 64.59 86.01 65.31 ;
      RECT 85.09 52.58 85.85 52.86 ;
      RECT 85.69 51.64 85.85 52.86 ;
      RECT 85.09 52.18 85.25 52.86 ;
      RECT 85.49 34.44 85.83 34.72 ;
      RECT 85.49 32.44 85.65 34.72 ;
      RECT 85.49 33.11 85.83 33.39 ;
      RECT 85.49 32.44 85.83 32.72 ;
      RECT 85.49 40.7 85.83 40.98 ;
      RECT 85.49 38.7 85.65 40.98 ;
      RECT 85.49 40.03 85.83 40.31 ;
      RECT 85.49 38.7 85.83 38.98 ;
      RECT 85.55 53.23 85.83 53.51 ;
      RECT 85.55 53.03 85.71 53.51 ;
      RECT 84.73 53.03 85.71 53.19 ;
      RECT 84.73 50.98 84.89 53.19 ;
      RECT 84.69 52.54 84.89 52.82 ;
      RECT 84.35 50.98 84.89 51.14 ;
      RECT 84.35 50.8 84.57 51.14 ;
      RECT 84.25 56.67 84.41 61.86 ;
      RECT 84.25 56.67 85.69 56.83 ;
      RECT 85.53 56 85.69 56.83 ;
      RECT 84.41 54.4 84.57 56.83 ;
      RECT 77.69 12.95 85.53 13.55 ;
      RECT 84.93 8.34 85.53 13.55 ;
      RECT 77.69 8.34 78.29 13.55 ;
      RECT 77.69 8.34 85.53 8.88 ;
      RECT 77.69 26.87 85.53 27.47 ;
      RECT 84.93 18.71 85.53 27.47 ;
      RECT 77.69 18.71 78.29 27.47 ;
      RECT 77.69 24.41 85.53 25.01 ;
      RECT 77.69 18.71 85.53 19.31 ;
      RECT 85.37 50.66 85.53 51.5 ;
      RECT 84.73 50.66 85.53 50.82 ;
      RECT 84.73 50.18 84.89 50.82 ;
      RECT 84.25 50.18 84.89 50.5 ;
      RECT 84.25 47.07 84.41 50.5 ;
      RECT 84.25 47.07 84.73 47.23 ;
      RECT 84.57 45.44 84.73 47.23 ;
      RECT 85.13 55.68 85.29 56.51 ;
      RECT 85.13 55.68 85.53 55.84 ;
      RECT 85.37 53.67 85.53 55.84 ;
      RECT 84.89 53.67 85.53 53.83 ;
      RECT 84.89 53.35 85.17 53.83 ;
      RECT 85.37 62.9 85.53 67.89 ;
      RECT 85.31 65.82 85.53 66.55 ;
      RECT 85.05 51.7 85.43 51.92 ;
      RECT 85.05 50.98 85.21 51.92 ;
      RECT 84.57 47.39 84.73 49.72 ;
      RECT 84.57 47.39 85.05 47.55 ;
      RECT 84.89 43.85 85.05 47.55 ;
      RECT 84.27 43.85 85.05 44.01 ;
      RECT 84.27 39.56 84.43 44.01 ;
      RECT 84.27 39.56 84.61 39.84 ;
      RECT 84.45 39.16 84.61 39.84 ;
      RECT 84.59 34.44 84.93 34.72 ;
      RECT 84.77 32.44 84.93 34.72 ;
      RECT 84.59 33.11 84.93 33.39 ;
      RECT 84.59 32.44 84.93 32.72 ;
      RECT 84.59 40.7 84.93 40.98 ;
      RECT 84.77 38.7 84.93 40.98 ;
      RECT 84.59 40.03 84.93 40.31 ;
      RECT 84.59 38.7 84.93 38.98 ;
      RECT 84.73 54.06 84.89 56.51 ;
      RECT 84.37 54.06 84.89 54.22 ;
      RECT 84.37 52.98 84.57 54.22 ;
      RECT 84.37 51.34 84.53 54.22 ;
      RECT 84.37 51.34 84.57 52.12 ;
      RECT 83.93 46.75 84.09 47.43 ;
      RECT 83.61 46.75 84.41 46.91 ;
      RECT 84.25 44.23 84.41 46.91 ;
      RECT 83.61 44.23 83.77 46.91 ;
      RECT 81.71 34.88 83.91 35.04 ;
      RECT 83.63 34.59 83.91 35.04 ;
      RECT 82.69 34.59 82.93 35.04 ;
      RECT 81.71 34.59 81.99 35.04 ;
      RECT 82.69 38.38 82.93 39.02 ;
      RECT 83.63 38.38 83.91 38.83 ;
      RECT 81.71 38.38 81.99 38.83 ;
      RECT 81.71 38.38 83.91 38.54 ;
      RECT 81.87 36.47 83.75 36.63 ;
      RECT 83.59 35.86 83.75 36.63 ;
      RECT 82.73 35.23 82.89 36.63 ;
      RECT 81.87 35.86 82.03 36.63 ;
      RECT 83.69 35.23 83.85 36.05 ;
      RECT 81.77 35.23 81.93 36.05 ;
      RECT 83.69 37.11 83.85 38.19 ;
      RECT 82.73 36.79 82.89 38.19 ;
      RECT 81.77 37.11 81.93 38.19 ;
      RECT 83.59 36.79 83.75 37.39 ;
      RECT 81.87 36.79 82.03 37.39 ;
      RECT 81.87 36.79 83.75 36.95 ;
      RECT 82.49 50.66 82.65 51.5 ;
      RECT 82.49 50.66 83.29 50.82 ;
      RECT 83.13 50.18 83.29 50.82 ;
      RECT 83.13 50.18 83.77 50.5 ;
      RECT 83.61 47.07 83.77 50.5 ;
      RECT 83.29 47.07 83.77 47.23 ;
      RECT 83.29 45.44 83.45 47.23 ;
      RECT 83.61 56.67 83.77 61.86 ;
      RECT 82.33 56.67 83.77 56.83 ;
      RECT 83.45 54.4 83.61 56.83 ;
      RECT 82.33 56 82.49 56.83 ;
      RECT 83.29 47.39 83.45 49.72 ;
      RECT 82.97 47.39 83.45 47.55 ;
      RECT 82.97 43.85 83.13 47.55 ;
      RECT 82.97 43.85 83.75 44.01 ;
      RECT 83.59 39.56 83.75 44.01 ;
      RECT 83.41 39.56 83.75 39.84 ;
      RECT 83.41 39.16 83.57 39.84 ;
      RECT 82.19 53.23 82.47 53.51 ;
      RECT 82.31 53.03 82.47 53.51 ;
      RECT 82.31 53.03 83.29 53.19 ;
      RECT 83.13 50.98 83.29 53.19 ;
      RECT 83.13 52.54 83.33 52.82 ;
      RECT 83.13 50.98 83.67 51.14 ;
      RECT 83.45 50.8 83.67 51.14 ;
      RECT 81.85 68.07 83.67 68.23 ;
      RECT 83.51 62.02 83.67 68.23 ;
      RECT 83.29 62.02 83.67 62.18 ;
      RECT 83.29 57.45 83.45 62.18 ;
      RECT 81.85 57.45 83.45 57.61 ;
      RECT 81.85 57.39 82.17 57.61 ;
      RECT 82.01 53.74 82.17 57.61 ;
      RECT 81.85 51.32 82.01 53.9 ;
      RECT 81.85 51.32 82.33 51.48 ;
      RECT 82.17 49.88 82.33 51.48 ;
      RECT 82.17 49.88 82.65 50.04 ;
      RECT 82.49 47.71 82.65 50.04 ;
      RECT 82.49 47.71 83.11 47.99 ;
      RECT 83.13 54.06 83.29 56.51 ;
      RECT 83.13 54.06 83.65 54.22 ;
      RECT 83.49 51.34 83.65 54.22 ;
      RECT 83.45 52.98 83.65 54.22 ;
      RECT 83.45 51.34 83.65 52.12 ;
      RECT 83.09 34.44 83.43 34.72 ;
      RECT 83.09 32.44 83.25 34.72 ;
      RECT 83.09 33.11 83.43 33.39 ;
      RECT 83.09 32.44 83.43 32.72 ;
      RECT 83.09 40.7 83.43 40.98 ;
      RECT 83.09 38.7 83.25 40.98 ;
      RECT 83.09 40.03 83.43 40.31 ;
      RECT 83.09 38.7 83.43 38.98 ;
      RECT 82.73 55.68 82.89 56.51 ;
      RECT 82.49 55.68 82.89 55.84 ;
      RECT 82.49 53.67 82.65 55.84 ;
      RECT 82.49 53.67 83.13 53.83 ;
      RECT 82.85 53.35 83.13 53.83 ;
      RECT 82.59 51.7 82.97 51.92 ;
      RECT 82.81 50.98 82.97 51.92 ;
      RECT 82.17 52.58 82.93 52.86 ;
      RECT 82.77 52.18 82.93 52.86 ;
      RECT 82.17 51.64 82.33 52.86 ;
      RECT 82.49 62.9 82.65 67.89 ;
      RECT 82.49 65.82 82.71 66.55 ;
      RECT 82.17 47.39 82.33 49.72 ;
      RECT 82.17 47.39 82.65 47.55 ;
      RECT 82.49 43.85 82.65 47.55 ;
      RECT 81.87 43.85 82.65 44.01 ;
      RECT 81.87 39.56 82.03 44.01 ;
      RECT 81.87 39.56 82.21 39.84 ;
      RECT 82.05 39.16 82.21 39.84 ;
      RECT 82.19 34.44 82.53 34.72 ;
      RECT 82.37 32.44 82.53 34.72 ;
      RECT 82.19 33.11 82.53 33.39 ;
      RECT 82.19 32.44 82.53 32.72 ;
      RECT 82.19 40.7 82.53 40.98 ;
      RECT 82.37 38.7 82.53 40.98 ;
      RECT 82.19 40.03 82.53 40.31 ;
      RECT 82.19 38.7 82.53 38.98 ;
      RECT 82.01 62.9 82.17 67.89 ;
      RECT 82.01 64.59 82.29 65.31 ;
      RECT 81.53 46.75 81.69 47.43 ;
      RECT 81.21 46.75 82.01 46.91 ;
      RECT 81.85 44.23 82.01 46.91 ;
      RECT 81.21 44.23 81.37 46.91 ;
      RECT 79.31 34.88 81.51 35.04 ;
      RECT 81.23 34.59 81.51 35.04 ;
      RECT 80.29 34.59 80.53 35.04 ;
      RECT 79.31 34.59 79.59 35.04 ;
      RECT 80.29 38.38 80.53 39.02 ;
      RECT 81.23 38.38 81.51 38.83 ;
      RECT 79.31 38.38 79.59 38.83 ;
      RECT 79.31 38.38 81.51 38.54 ;
      RECT 79.47 36.47 81.35 36.63 ;
      RECT 81.19 35.88 81.35 36.63 ;
      RECT 80.33 35.23 80.49 36.63 ;
      RECT 79.47 35.88 79.63 36.63 ;
      RECT 81.29 35.23 81.45 36.06 ;
      RECT 79.37 35.23 79.53 36.06 ;
      RECT 81.29 37.11 81.45 38.19 ;
      RECT 80.33 36.79 80.49 38.19 ;
      RECT 79.37 37.11 79.53 38.19 ;
      RECT 81.19 36.79 81.35 37.39 ;
      RECT 79.47 36.79 79.63 37.39 ;
      RECT 79.47 36.79 81.35 36.95 ;
      RECT 79.55 68.07 81.37 68.23 ;
      RECT 79.55 62.02 79.71 68.23 ;
      RECT 79.55 62.02 79.93 62.18 ;
      RECT 79.77 57.45 79.93 62.18 ;
      RECT 79.77 57.45 81.37 57.61 ;
      RECT 81.05 57.39 81.37 57.61 ;
      RECT 81.05 53.74 81.21 57.61 ;
      RECT 81.21 51.32 81.37 53.9 ;
      RECT 80.89 51.32 81.37 51.48 ;
      RECT 80.89 49.88 81.05 51.48 ;
      RECT 80.57 49.88 81.05 50.04 ;
      RECT 80.57 47.71 80.73 50.04 ;
      RECT 80.11 47.71 80.73 47.99 ;
      RECT 80.89 47.39 81.05 49.72 ;
      RECT 80.57 47.39 81.05 47.55 ;
      RECT 80.57 43.85 80.73 47.55 ;
      RECT 80.57 43.85 81.35 44.01 ;
      RECT 81.19 39.56 81.35 44.01 ;
      RECT 81.01 39.56 81.35 39.84 ;
      RECT 81.01 39.16 81.17 39.84 ;
      RECT 81.05 62.9 81.21 67.89 ;
      RECT 80.93 64.59 81.21 65.31 ;
      RECT 80.29 52.58 81.05 52.86 ;
      RECT 80.89 51.64 81.05 52.86 ;
      RECT 80.29 52.18 80.45 52.86 ;
      RECT 80.69 34.44 81.03 34.72 ;
      RECT 80.69 32.44 80.85 34.72 ;
      RECT 80.69 33.11 81.03 33.39 ;
      RECT 80.69 32.44 81.03 32.72 ;
      RECT 80.69 40.7 81.03 40.98 ;
      RECT 80.69 38.7 80.85 40.98 ;
      RECT 80.69 40.03 81.03 40.31 ;
      RECT 80.69 38.7 81.03 38.98 ;
      RECT 80.75 53.23 81.03 53.51 ;
      RECT 80.75 53.03 80.91 53.51 ;
      RECT 79.93 53.03 80.91 53.19 ;
      RECT 79.93 50.98 80.09 53.19 ;
      RECT 79.89 52.54 80.09 52.82 ;
      RECT 79.55 50.98 80.09 51.14 ;
      RECT 79.55 50.8 79.77 51.14 ;
      RECT 79.45 56.67 79.61 61.86 ;
      RECT 79.45 56.67 80.89 56.83 ;
      RECT 80.73 56 80.89 56.83 ;
      RECT 79.61 54.4 79.77 56.83 ;
      RECT 80.57 50.66 80.73 51.5 ;
      RECT 79.93 50.66 80.73 50.82 ;
      RECT 79.93 50.18 80.09 50.82 ;
      RECT 79.45 50.18 80.09 50.5 ;
      RECT 79.45 47.07 79.61 50.5 ;
      RECT 79.45 47.07 79.93 47.23 ;
      RECT 79.77 45.44 79.93 47.23 ;
      RECT 80.33 55.68 80.49 56.51 ;
      RECT 80.33 55.68 80.73 55.84 ;
      RECT 80.57 53.67 80.73 55.84 ;
      RECT 80.09 53.67 80.73 53.83 ;
      RECT 80.09 53.35 80.37 53.83 ;
      RECT 80.57 62.9 80.73 67.89 ;
      RECT 80.51 65.82 80.73 66.55 ;
      RECT 80.25 51.7 80.63 51.92 ;
      RECT 80.25 50.98 80.41 51.92 ;
      RECT 79.77 47.39 79.93 49.72 ;
      RECT 79.77 47.39 80.25 47.55 ;
      RECT 80.09 43.85 80.25 47.55 ;
      RECT 79.47 43.85 80.25 44.01 ;
      RECT 79.47 39.56 79.63 44.01 ;
      RECT 79.47 39.56 79.81 39.84 ;
      RECT 79.65 39.16 79.81 39.84 ;
      RECT 79.79 34.44 80.13 34.72 ;
      RECT 79.97 32.44 80.13 34.72 ;
      RECT 79.79 33.11 80.13 33.39 ;
      RECT 79.79 32.44 80.13 32.72 ;
      RECT 79.79 40.7 80.13 40.98 ;
      RECT 79.97 38.7 80.13 40.98 ;
      RECT 79.79 40.03 80.13 40.31 ;
      RECT 79.79 38.7 80.13 38.98 ;
      RECT 79.93 54.06 80.09 56.51 ;
      RECT 79.57 54.06 80.09 54.22 ;
      RECT 79.57 52.98 79.77 54.22 ;
      RECT 79.57 51.34 79.73 54.22 ;
      RECT 79.57 51.34 79.77 52.12 ;
      RECT 79.13 46.75 79.29 47.43 ;
      RECT 78.81 46.75 79.61 46.91 ;
      RECT 79.45 44.23 79.61 46.91 ;
      RECT 78.81 44.23 78.97 46.91 ;
      RECT 76.91 34.88 79.11 35.04 ;
      RECT 78.83 34.59 79.11 35.04 ;
      RECT 77.89 34.59 78.13 35.04 ;
      RECT 76.91 34.59 77.19 35.04 ;
      RECT 77.89 38.38 78.13 39.02 ;
      RECT 78.83 38.38 79.11 38.83 ;
      RECT 76.91 38.38 77.19 38.83 ;
      RECT 76.91 38.38 79.11 38.54 ;
      RECT 77.07 36.47 78.95 36.63 ;
      RECT 78.79 35.86 78.95 36.63 ;
      RECT 77.93 35.23 78.09 36.63 ;
      RECT 77.07 35.86 77.23 36.63 ;
      RECT 78.89 35.23 79.05 36.05 ;
      RECT 76.97 35.23 77.13 36.05 ;
      RECT 78.89 37.11 79.05 38.19 ;
      RECT 77.93 36.79 78.09 38.19 ;
      RECT 76.97 37.11 77.13 38.19 ;
      RECT 78.79 36.79 78.95 37.39 ;
      RECT 77.07 36.79 77.23 37.39 ;
      RECT 77.07 36.79 78.95 36.95 ;
      RECT 77.69 50.66 77.85 51.5 ;
      RECT 77.69 50.66 78.49 50.82 ;
      RECT 78.33 50.18 78.49 50.82 ;
      RECT 78.33 50.18 78.97 50.5 ;
      RECT 78.81 47.07 78.97 50.5 ;
      RECT 78.49 47.07 78.97 47.23 ;
      RECT 78.49 45.44 78.65 47.23 ;
      RECT 78.81 56.67 78.97 61.86 ;
      RECT 77.53 56.67 78.97 56.83 ;
      RECT 78.65 54.4 78.81 56.83 ;
      RECT 77.53 56 77.69 56.83 ;
      RECT 78.49 47.39 78.65 49.72 ;
      RECT 78.17 47.39 78.65 47.55 ;
      RECT 78.17 43.85 78.33 47.55 ;
      RECT 78.17 43.85 78.95 44.01 ;
      RECT 78.79 39.56 78.95 44.01 ;
      RECT 78.61 39.56 78.95 39.84 ;
      RECT 78.61 39.16 78.77 39.84 ;
      RECT 77.39 53.23 77.67 53.51 ;
      RECT 77.51 53.03 77.67 53.51 ;
      RECT 77.51 53.03 78.49 53.19 ;
      RECT 78.33 50.98 78.49 53.19 ;
      RECT 78.33 52.54 78.53 52.82 ;
      RECT 78.33 50.98 78.87 51.14 ;
      RECT 78.65 50.8 78.87 51.14 ;
      RECT 77.05 68.07 78.87 68.23 ;
      RECT 78.71 62.02 78.87 68.23 ;
      RECT 78.49 62.02 78.87 62.18 ;
      RECT 78.49 57.45 78.65 62.18 ;
      RECT 77.05 57.45 78.65 57.61 ;
      RECT 77.05 57.39 77.37 57.61 ;
      RECT 77.21 53.74 77.37 57.61 ;
      RECT 77.05 51.32 77.21 53.9 ;
      RECT 77.05 51.32 77.53 51.48 ;
      RECT 77.37 49.88 77.53 51.48 ;
      RECT 77.37 49.88 77.85 50.04 ;
      RECT 77.69 47.71 77.85 50.04 ;
      RECT 77.69 47.71 78.31 47.99 ;
      RECT 78.33 54.06 78.49 56.51 ;
      RECT 78.33 54.06 78.85 54.22 ;
      RECT 78.69 51.34 78.85 54.22 ;
      RECT 78.65 52.98 78.85 54.22 ;
      RECT 78.65 51.34 78.85 52.12 ;
      RECT 78.29 34.44 78.63 34.72 ;
      RECT 78.29 32.44 78.45 34.72 ;
      RECT 78.29 33.11 78.63 33.39 ;
      RECT 78.29 32.44 78.63 32.72 ;
      RECT 78.29 40.7 78.63 40.98 ;
      RECT 78.29 38.7 78.45 40.98 ;
      RECT 78.29 40.03 78.63 40.31 ;
      RECT 78.29 38.7 78.63 38.98 ;
      RECT 77.93 55.68 78.09 56.51 ;
      RECT 77.69 55.68 78.09 55.84 ;
      RECT 77.69 53.67 77.85 55.84 ;
      RECT 77.69 53.67 78.33 53.83 ;
      RECT 78.05 53.35 78.33 53.83 ;
      RECT 77.79 51.7 78.17 51.92 ;
      RECT 78.01 50.98 78.17 51.92 ;
      RECT 77.37 52.58 78.13 52.86 ;
      RECT 77.97 52.18 78.13 52.86 ;
      RECT 77.37 51.64 77.53 52.86 ;
      RECT 77.69 62.9 77.85 67.89 ;
      RECT 77.69 65.82 77.91 66.55 ;
      RECT 77.37 47.39 77.53 49.72 ;
      RECT 77.37 47.39 77.85 47.55 ;
      RECT 77.69 43.85 77.85 47.55 ;
      RECT 77.07 43.85 77.85 44.01 ;
      RECT 77.07 39.56 77.23 44.01 ;
      RECT 77.07 39.56 77.41 39.84 ;
      RECT 77.25 39.16 77.41 39.84 ;
      RECT 77.39 34.44 77.73 34.72 ;
      RECT 77.57 32.44 77.73 34.72 ;
      RECT 77.39 33.11 77.73 33.39 ;
      RECT 77.39 32.44 77.73 32.72 ;
      RECT 77.39 40.7 77.73 40.98 ;
      RECT 77.57 38.7 77.73 40.98 ;
      RECT 77.39 40.03 77.73 40.31 ;
      RECT 77.39 38.7 77.73 38.98 ;
      RECT 77.21 62.9 77.37 67.89 ;
      RECT 77.21 64.59 77.49 65.31 ;
      RECT 76.73 46.75 76.89 47.43 ;
      RECT 76.41 46.75 77.21 46.91 ;
      RECT 77.05 44.23 77.21 46.91 ;
      RECT 76.41 44.23 76.57 46.91 ;
      RECT 76.21 10.08 76.37 11.89 ;
      RECT 76.21 10.08 76.95 10.24 ;
      RECT 76.73 8.88 76.89 10.24 ;
      RECT 76.73 7.5 76.89 8.72 ;
      RECT 76.68 7.58 76.89 7.9 ;
      RECT 75.65 7.59 76.89 7.75 ;
      RECT 76.61 7.58 76.89 7.75 ;
      RECT 68.69 15.8 68.85 16.08 ;
      RECT 65.57 15.8 65.73 16.08 ;
      RECT 68.09 15.8 68.85 15.96 ;
      RECT 65.57 15.8 66.33 15.96 ;
      RECT 66.17 14.07 66.33 15.96 ;
      RECT 74.59 14.25 74.75 15.89 ;
      RECT 59.67 14.25 59.83 15.89 ;
      RECT 67.13 12.21 67.29 15.8 ;
      RECT 68.09 14.07 68.25 15.96 ;
      RECT 72.07 14.12 72.25 15.79 ;
      RECT 70.79 14.1 70.95 15.79 ;
      RECT 63.47 14.1 63.63 15.79 ;
      RECT 62.17 14.12 62.35 15.79 ;
      RECT 75.93 14.64 76.09 15.6 ;
      RECT 58.33 14.64 58.49 15.6 ;
      RECT 76.73 12.64 76.89 14.96 ;
      RECT 57.53 12.64 57.69 14.96 ;
      RECT 69.75 14.1 69.91 14.89 ;
      RECT 64.51 14.1 64.67 14.89 ;
      RECT 74.31 14.64 76.89 14.84 ;
      RECT 57.53 14.64 60.11 14.84 ;
      RECT 59.95 12.56 60.11 14.84 ;
      RECT 74.31 14.25 75.76 14.84 ;
      RECT 58.66 14.25 60.11 14.84 ;
      RECT 68.81 14.36 69.91 14.52 ;
      RECT 64.51 14.36 65.61 14.52 ;
      RECT 65.45 14.08 65.61 14.52 ;
      RECT 68.81 14.08 68.97 14.52 ;
      RECT 70.79 14.12 74.47 14.28 ;
      RECT 58.66 14.25 63.63 14.28 ;
      RECT 69.75 14.1 71.27 14.26 ;
      RECT 63.15 14.1 64.67 14.26 ;
      RECT 59.95 14.12 64.67 14.26 ;
      RECT 68.09 14.08 68.97 14.24 ;
      RECT 65.45 14.08 66.33 14.24 ;
      RECT 65.99 14.07 68.43 14.23 ;
      RECT 74.31 12.56 74.47 14.84 ;
      RECT 73.35 12.55 73.51 14.28 ;
      RECT 72.47 13.45 72.63 14.28 ;
      RECT 61.79 13.45 61.95 14.28 ;
      RECT 60.91 12.55 61.07 14.28 ;
      RECT 70.01 12.32 70.17 14.26 ;
      RECT 64.25 12.32 64.41 14.26 ;
      RECT 68.27 13.38 68.43 14.24 ;
      RECT 65.99 13.38 66.15 14.24 ;
      RECT 72.39 12.55 72.55 13.61 ;
      RECT 61.87 12.55 62.03 13.61 ;
      RECT 68.15 13.38 68.43 13.54 ;
      RECT 65.99 13.38 66.27 13.54 ;
      RECT 76.06 17.18 76.22 18.9 ;
      RECT 76.06 17.96 76.89 18.12 ;
      RECT 76.73 17.84 76.89 18.12 ;
      RECT 76.02 17.06 76.18 17.34 ;
      RECT 75.04 19.61 75.2 21.25 ;
      RECT 68.09 20.42 68.25 21.25 ;
      RECT 67.13 16.39 67.29 21.25 ;
      RECT 66.17 20.42 66.33 21.25 ;
      RECT 59.22 19.61 59.38 21.25 ;
      RECT 75.82 20.89 76.24 21.05 ;
      RECT 74.08 19.61 74.24 21.05 ;
      RECT 60.18 19.61 60.34 21.05 ;
      RECT 58.18 20.89 58.6 21.05 ;
      RECT 58.44 19.61 58.6 21.05 ;
      RECT 73.08 20.21 73.24 20.89 ;
      RECT 70.83 20.43 70.99 20.89 ;
      RECT 63.43 20.43 63.59 20.89 ;
      RECT 61.18 20.21 61.34 20.89 ;
      RECT 75.82 19.61 75.98 21.05 ;
      RECT 70.37 20.43 70.99 20.59 ;
      RECT 63.43 20.43 64.05 20.59 ;
      RECT 63.89 19.1 64.05 20.59 ;
      RECT 68.17 19.16 68.33 20.58 ;
      RECT 66.09 19.16 66.25 20.58 ;
      RECT 69.41 19.16 69.57 20.49 ;
      RECT 64.85 19.16 65.01 20.49 ;
      RECT 70.37 19.1 70.53 20.59 ;
      RECT 73.08 20.21 74.24 20.37 ;
      RECT 74.04 19.61 74.24 20.37 ;
      RECT 60.18 20.21 61.34 20.37 ;
      RECT 60.18 19.61 60.38 20.37 ;
      RECT 74.04 19.61 75.2 19.81 ;
      RECT 59.22 19.61 60.38 19.81 ;
      RECT 73.87 19.61 76.81 19.77 ;
      RECT 57.61 19.61 60.55 19.77 ;
      RECT 60.39 19.1 60.55 19.77 ;
      RECT 72.91 19.1 73.19 19.73 ;
      RECT 61.23 19.1 61.51 19.73 ;
      RECT 73.87 19.1 74.03 19.77 ;
      RECT 69.41 19.16 70.53 19.37 ;
      RECT 63.89 19.16 65.01 19.37 ;
      RECT 63.89 19.16 70.53 19.32 ;
      RECT 69.52 19.1 74.03 19.26 ;
      RECT 69.05 18.46 69.21 19.32 ;
      RECT 68.09 17.56 68.25 19.32 ;
      RECT 66.17 17.56 66.33 19.32 ;
      RECT 65.21 18.46 65.37 19.32 ;
      RECT 60.39 19.1 64.9 19.26 ;
      RECT 63.76 17.76 63.92 19.26 ;
      RECT 70.5 19.01 72.42 19.26 ;
      RECT 72.24 16.65 72.42 19.26 ;
      RECT 62 19.01 63.92 19.26 ;
      RECT 71.3 17.58 71.46 19.26 ;
      RECT 70.5 17.76 70.66 19.26 ;
      RECT 62.96 17.58 63.12 19.26 ;
      RECT 62 16.65 62.18 19.26 ;
      RECT 69.97 17.76 70.66 17.92 ;
      RECT 63.76 17.76 64.45 17.92 ;
      RECT 64.29 16.77 64.45 17.92 ;
      RECT 69.97 16.77 70.13 17.92 ;
      RECT 76.5 15.57 76.66 17.28 ;
      RECT 75.9 16.43 76.06 16.71 ;
      RECT 75.9 16.43 76.66 16.59 ;
      RECT 76.44 15.57 76.72 15.73 ;
      RECT 74.51 34.88 76.71 35.04 ;
      RECT 76.43 34.59 76.71 35.04 ;
      RECT 75.49 34.59 75.73 35.04 ;
      RECT 74.51 34.59 74.79 35.04 ;
      RECT 75.49 38.38 75.73 39.02 ;
      RECT 76.43 38.38 76.71 38.83 ;
      RECT 74.51 38.38 74.79 38.83 ;
      RECT 74.51 38.38 76.71 38.54 ;
      RECT 76.03 23.66 76.57 23.82 ;
      RECT 76.41 20.12 76.57 23.82 ;
      RECT 76.11 23.22 76.57 23.38 ;
      RECT 76.41 20.83 76.66 21.11 ;
      RECT 76.14 20.12 76.57 20.28 ;
      RECT 76.46 26.15 76.62 28.96 ;
      RECT 76.46 26.15 76.65 26.51 ;
      RECT 74.67 36.47 76.55 36.63 ;
      RECT 76.39 35.88 76.55 36.63 ;
      RECT 75.53 35.23 75.69 36.63 ;
      RECT 74.67 35.88 74.83 36.63 ;
      RECT 76.49 35.23 76.65 36.06 ;
      RECT 74.57 35.23 74.73 36.06 ;
      RECT 76.49 37.11 76.65 38.19 ;
      RECT 75.53 36.79 75.69 38.19 ;
      RECT 74.57 37.11 74.73 38.19 ;
      RECT 76.39 36.79 76.55 37.39 ;
      RECT 74.67 36.79 74.83 37.39 ;
      RECT 74.67 36.79 76.55 36.95 ;
      RECT 74.75 68.07 76.57 68.23 ;
      RECT 74.75 62.02 74.91 68.23 ;
      RECT 74.75 62.02 75.13 62.18 ;
      RECT 74.97 57.45 75.13 62.18 ;
      RECT 74.97 57.45 76.57 57.61 ;
      RECT 76.25 57.39 76.57 57.61 ;
      RECT 76.25 53.74 76.41 57.61 ;
      RECT 76.41 51.32 76.57 53.9 ;
      RECT 76.09 51.32 76.57 51.48 ;
      RECT 76.09 49.88 76.25 51.48 ;
      RECT 75.77 49.88 76.25 50.04 ;
      RECT 75.77 47.71 75.93 50.04 ;
      RECT 75.31 47.71 75.93 47.99 ;
      RECT 76.09 47.39 76.25 49.72 ;
      RECT 75.77 47.39 76.25 47.55 ;
      RECT 75.77 43.85 75.93 47.55 ;
      RECT 75.77 43.85 76.55 44.01 ;
      RECT 76.39 39.56 76.55 44.01 ;
      RECT 76.21 39.56 76.55 39.84 ;
      RECT 76.21 39.16 76.37 39.84 ;
      RECT 73.91 8.96 74.23 9.12 ;
      RECT 73.91 7.8 74.07 9.12 ;
      RECT 76.25 7.91 76.41 8.8 ;
      RECT 75.33 7.91 76.41 8.07 ;
      RECT 73.91 7.8 75.49 7.96 ;
      RECT 76.23 23.98 76.41 24.52 ;
      RECT 75.71 23.98 76.41 24.14 ;
      RECT 75.71 23.27 75.87 24.14 ;
      RECT 75.77 21.78 75.93 23.43 ;
      RECT 75.63 21.21 75.79 21.94 ;
      RECT 75.5 20.95 75.66 21.37 ;
      RECT 76.25 62.9 76.41 67.89 ;
      RECT 76.13 64.59 76.41 65.31 ;
      RECT 75.49 52.58 76.25 52.86 ;
      RECT 76.09 51.64 76.25 52.86 ;
      RECT 75.49 52.18 75.65 52.86 ;
      RECT 75.89 34.44 76.23 34.72 ;
      RECT 75.89 32.44 76.05 34.72 ;
      RECT 75.89 33.11 76.23 33.39 ;
      RECT 75.89 32.44 76.23 32.72 ;
      RECT 75.89 40.7 76.23 40.98 ;
      RECT 75.89 38.7 76.05 40.98 ;
      RECT 75.89 40.03 76.23 40.31 ;
      RECT 75.89 38.7 76.23 38.98 ;
      RECT 75.95 53.23 76.23 53.51 ;
      RECT 75.95 53.03 76.11 53.51 ;
      RECT 75.13 53.03 76.11 53.19 ;
      RECT 75.13 50.98 75.29 53.19 ;
      RECT 75.09 52.54 75.29 52.82 ;
      RECT 74.75 50.98 75.29 51.14 ;
      RECT 74.75 50.8 74.97 51.14 ;
      RECT 75.13 28.52 76.22 28.68 ;
      RECT 75.13 28.35 75.41 28.68 ;
      RECT 74.73 28.35 75.41 28.51 ;
      RECT 75.98 24.79 76.14 28.32 ;
      RECT 75.45 25.16 76.14 25.32 ;
      RECT 75.93 12.92 76.09 13.67 ;
      RECT 75.73 12.92 76.09 13.08 ;
      RECT 75.73 9.68 75.89 13.08 ;
      RECT 75.73 9.68 75.93 11.89 ;
      RECT 74.95 9.68 75.93 9.84 ;
      RECT 74.95 8.6 75.11 9.84 ;
      RECT 74.65 56.67 74.81 61.86 ;
      RECT 74.65 56.67 76.09 56.83 ;
      RECT 75.93 56 76.09 56.83 ;
      RECT 74.81 54.4 74.97 56.83 ;
      RECT 74.09 26.02 74.65 26.18 ;
      RECT 74.49 25.58 74.65 26.18 ;
      RECT 74.49 25.58 75.19 25.74 ;
      RECT 75.03 22.71 75.19 25.74 ;
      RECT 74.99 24 75.19 25.74 ;
      RECT 74.99 24.3 75.99 24.46 ;
      RECT 74.93 22.04 75.09 22.99 ;
      RECT 74.77 21.85 74.93 22.32 ;
      RECT 75.77 50.66 75.93 51.5 ;
      RECT 75.13 50.66 75.93 50.82 ;
      RECT 75.13 50.18 75.29 50.82 ;
      RECT 74.65 50.18 75.29 50.5 ;
      RECT 74.65 47.07 74.81 50.5 ;
      RECT 74.65 47.07 75.13 47.23 ;
      RECT 74.97 45.44 75.13 47.23 ;
      RECT 75.53 55.68 75.69 56.51 ;
      RECT 75.53 55.68 75.93 55.84 ;
      RECT 75.77 53.67 75.93 55.84 ;
      RECT 75.29 53.67 75.93 53.83 ;
      RECT 75.29 53.35 75.57 53.83 ;
      RECT 75.77 62.9 75.93 67.89 ;
      RECT 75.71 65.82 75.93 66.55 ;
      RECT 75.45 51.7 75.83 51.92 ;
      RECT 75.45 50.98 75.61 51.92 ;
      RECT 72.87 26.36 73.03 26.72 ;
      RECT 72.87 26.36 75.17 26.52 ;
      RECT 75.01 26.04 75.17 26.52 ;
      RECT 75.01 26.04 75.82 26.2 ;
      RECT 75.58 16.52 75.74 18.9 ;
      RECT 75.38 16.52 75.74 16.8 ;
      RECT 75.45 15.31 75.61 16.8 ;
      RECT 75.25 22.13 75.61 22.41 ;
      RECT 75.25 21.53 75.41 22.41 ;
      RECT 74.38 21.53 74.54 21.92 ;
      RECT 74.38 21.53 75.41 21.69 ;
      RECT 74.56 20.21 74.72 21.69 ;
      RECT 75.41 11.5 75.57 13.22 ;
      RECT 74.05 12.22 75.57 12.38 ;
      RECT 75.15 11.5 75.57 11.66 ;
      RECT 74.97 47.39 75.13 49.72 ;
      RECT 74.97 47.39 75.45 47.55 ;
      RECT 75.29 43.85 75.45 47.55 ;
      RECT 74.67 43.85 75.45 44.01 ;
      RECT 74.67 39.56 74.83 44.01 ;
      RECT 74.67 39.56 75.01 39.84 ;
      RECT 74.85 39.16 75.01 39.84 ;
      RECT 74.48 18.3 75.42 18.46 ;
      RECT 75.06 17.05 75.42 18.46 ;
      RECT 75.06 16.2 75.22 18.46 ;
      RECT 74.31 16.2 75.27 16.36 ;
      RECT 75.11 16.08 75.27 16.36 ;
      RECT 73.87 16.07 74.54 16.23 ;
      RECT 74.99 34.44 75.33 34.72 ;
      RECT 75.17 32.44 75.33 34.72 ;
      RECT 74.99 33.11 75.33 33.39 ;
      RECT 74.99 32.44 75.33 32.72 ;
      RECT 74.99 40.7 75.33 40.98 ;
      RECT 75.17 38.7 75.33 40.98 ;
      RECT 74.99 40.03 75.33 40.31 ;
      RECT 74.99 38.7 75.33 38.98 ;
      RECT 75.13 54.06 75.29 56.51 ;
      RECT 74.77 54.06 75.29 54.22 ;
      RECT 74.77 52.98 74.97 54.22 ;
      RECT 74.77 51.34 74.93 54.22 ;
      RECT 74.77 51.34 74.97 52.12 ;
      RECT 73.04 28.01 75.2 28.17 ;
      RECT 75.04 26.68 75.2 28.17 ;
      RECT 74.04 26.97 74.2 28.17 ;
      RECT 73.04 27.93 73.36 28.17 ;
      RECT 73.04 27.34 73.2 28.17 ;
      RECT 73.83 12.56 73.99 13.61 ;
      RECT 73.73 11.9 73.89 13.24 ;
      RECT 73.73 11.9 75.01 12.06 ;
      RECT 73.91 9.6 74.07 12.06 ;
      RECT 74.72 16.52 74.9 16.84 ;
      RECT 74 16.52 74.9 16.68 ;
      RECT 74.71 23.18 74.87 23.84 ;
      RECT 74.54 23.18 74.87 23.34 ;
      RECT 74.54 22.65 74.7 23.34 ;
      RECT 74.33 46.75 74.49 47.43 ;
      RECT 74.01 46.75 74.81 46.91 ;
      RECT 74.65 44.23 74.81 46.91 ;
      RECT 74.01 44.23 74.17 46.91 ;
      RECT 74.52 26.69 74.68 27.85 ;
      RECT 74.48 26.69 74.72 27.33 ;
      RECT 74.39 9.28 74.55 11.72 ;
      RECT 73.43 8.12 73.59 11.72 ;
      RECT 72.47 8.5 72.63 11.72 ;
      RECT 70.81 9.63 70.97 11.4 ;
      RECT 70.81 9.95 72.63 10.11 ;
      RECT 71.5 9.79 71.66 10.11 ;
      RECT 74.43 8.12 74.63 9.84 ;
      RECT 70.75 9.63 71.26 9.79 ;
      RECT 73.43 9.28 74.63 9.44 ;
      RECT 72.43 8.5 72.74 8.78 ;
      RECT 72.43 8.56 73.59 8.72 ;
      RECT 69.45 28.74 74.57 28.9 ;
      RECT 72.65 27.92 72.81 28.9 ;
      RECT 71.21 27.92 71.37 28.9 ;
      RECT 74.26 16.92 74.42 18.12 ;
      RECT 74.02 16.92 74.42 17.08 ;
      RECT 72.11 34.88 74.31 35.04 ;
      RECT 74.03 34.59 74.31 35.04 ;
      RECT 73.09 34.59 73.33 35.04 ;
      RECT 72.11 34.59 72.39 35.04 ;
      RECT 73.09 38.38 73.33 39.02 ;
      RECT 74.03 38.38 74.31 38.83 ;
      RECT 72.11 38.38 72.39 38.83 ;
      RECT 72.11 38.38 74.31 38.54 ;
      RECT 71.93 21.69 72.09 26.21 ;
      RECT 73.17 24.34 73.33 26.2 ;
      RECT 70.69 24.35 70.85 26.2 ;
      RECT 74.05 24.04 74.27 25.52 ;
      RECT 69.75 24.04 69.97 25.52 ;
      RECT 73.17 24.46 74.27 24.63 ;
      RECT 69.75 24.46 70.85 24.63 ;
      RECT 70.67 21.69 70.83 24.63 ;
      RECT 73.19 21.69 73.35 24.63 ;
      RECT 70.67 21.69 73.35 21.85 ;
      RECT 72.27 36.47 74.15 36.63 ;
      RECT 73.99 35.86 74.15 36.63 ;
      RECT 73.13 35.23 73.29 36.63 ;
      RECT 72.27 35.86 72.43 36.63 ;
      RECT 74.09 35.23 74.25 36.05 ;
      RECT 72.17 35.23 72.33 36.05 ;
      RECT 74.09 37.11 74.25 38.19 ;
      RECT 73.13 36.79 73.29 38.19 ;
      RECT 72.17 37.11 72.33 38.19 ;
      RECT 73.99 36.79 74.15 37.39 ;
      RECT 72.27 36.79 72.43 37.39 ;
      RECT 72.27 36.79 74.15 36.95 ;
      RECT 74.05 21.37 74.21 23.37 ;
      RECT 70.21 21.37 74.21 21.53 ;
      RECT 73.56 20.73 73.72 21.53 ;
      RECT 70.21 20.78 70.37 21.53 ;
      RECT 72.89 50.66 73.05 51.5 ;
      RECT 72.89 50.66 73.69 50.82 ;
      RECT 73.53 50.18 73.69 50.82 ;
      RECT 73.53 50.18 74.17 50.5 ;
      RECT 74.01 47.07 74.17 50.5 ;
      RECT 73.69 47.07 74.17 47.23 ;
      RECT 73.69 45.44 73.85 47.23 ;
      RECT 74.01 56.67 74.17 61.86 ;
      RECT 72.73 56.67 74.17 56.83 ;
      RECT 73.85 54.4 74.01 56.83 ;
      RECT 72.73 56 72.89 56.83 ;
      RECT 73.69 47.39 73.85 49.72 ;
      RECT 73.37 47.39 73.85 47.55 ;
      RECT 73.37 43.85 73.53 47.55 ;
      RECT 73.37 43.85 74.15 44.01 ;
      RECT 73.99 39.56 74.15 44.01 ;
      RECT 73.81 39.56 74.15 39.84 ;
      RECT 73.81 39.16 73.97 39.84 ;
      RECT 72.59 53.23 72.87 53.51 ;
      RECT 72.71 53.03 72.87 53.51 ;
      RECT 72.71 53.03 73.69 53.19 ;
      RECT 73.53 50.98 73.69 53.19 ;
      RECT 73.53 52.54 73.73 52.82 ;
      RECT 73.53 50.98 74.07 51.14 ;
      RECT 73.85 50.8 74.07 51.14 ;
      RECT 72.25 68.07 74.07 68.23 ;
      RECT 73.91 62.02 74.07 68.23 ;
      RECT 73.69 62.02 74.07 62.18 ;
      RECT 73.69 57.45 73.85 62.18 ;
      RECT 72.25 57.45 73.85 57.61 ;
      RECT 72.25 57.39 72.57 57.61 ;
      RECT 72.41 53.74 72.57 57.61 ;
      RECT 72.25 51.32 72.41 53.9 ;
      RECT 72.25 51.32 72.73 51.48 ;
      RECT 72.57 49.88 72.73 51.48 ;
      RECT 72.57 49.88 73.05 50.04 ;
      RECT 72.89 47.71 73.05 50.04 ;
      RECT 72.89 47.71 73.51 47.99 ;
      RECT 73.53 54.06 73.69 56.51 ;
      RECT 73.53 54.06 74.05 54.22 ;
      RECT 73.89 51.34 74.05 54.22 ;
      RECT 73.85 52.98 74.05 54.22 ;
      RECT 73.85 51.34 74.05 52.12 ;
      RECT 72.74 18.78 73.86 18.94 ;
      RECT 73.68 17.48 73.86 18.94 ;
      RECT 71.78 17.26 71.95 18.8 ;
      RECT 71.79 16.12 71.95 18.8 ;
      RECT 70.82 16.44 70.98 18.8 ;
      RECT 72.74 16.03 72.9 18.94 ;
      RECT 70.77 16.44 70.98 17.57 ;
      RECT 73.68 16.44 73.84 18.94 ;
      RECT 70.77 17.26 71.95 17.42 ;
      RECT 70.77 16.44 71.05 17.42 ;
      RECT 73.55 14.52 73.71 16.71 ;
      RECT 69.77 16.12 72.9 16.28 ;
      RECT 72.59 14.52 72.75 16.28 ;
      RECT 71.59 14.84 71.75 16.28 ;
      RECT 72.59 14.52 73.71 14.68 ;
      RECT 73.49 34.44 73.83 34.72 ;
      RECT 73.49 32.44 73.65 34.72 ;
      RECT 73.49 33.11 73.83 33.39 ;
      RECT 73.49 32.44 73.83 32.72 ;
      RECT 73.49 40.7 73.83 40.98 ;
      RECT 73.49 38.7 73.65 40.98 ;
      RECT 73.49 40.03 73.83 40.31 ;
      RECT 73.49 38.7 73.83 38.98 ;
      RECT 73.65 21.85 73.81 24.3 ;
      RECT 73.51 21.85 73.81 22.13 ;
      RECT 73.49 24.79 73.69 25.35 ;
      RECT 73.49 24.79 73.81 25.03 ;
      RECT 72.17 28.04 72.49 28.32 ;
      RECT 72.33 25.99 72.49 28.32 ;
      RECT 73.52 27.02 73.68 27.7 ;
      RECT 72.33 27.02 73.68 27.18 ;
      RECT 72.33 25.99 72.71 26.23 ;
      RECT 72.55 25.16 72.71 26.23 ;
      RECT 72.19 20.26 72.35 21.05 ;
      RECT 72.19 20.26 72.92 20.44 ;
      RECT 72.76 19.89 72.92 20.44 ;
      RECT 72.76 19.89 73.58 20.05 ;
      RECT 73.39 19.61 73.58 20.05 ;
      RECT 73.39 19.61 73.67 19.77 ;
      RECT 73.13 55.68 73.29 56.51 ;
      RECT 72.89 55.68 73.29 55.84 ;
      RECT 72.89 53.67 73.05 55.84 ;
      RECT 72.89 53.67 73.53 53.83 ;
      RECT 73.25 53.35 73.53 53.83 ;
      RECT 72.99 51.7 73.37 51.92 ;
      RECT 73.21 50.98 73.37 51.92 ;
      RECT 72.57 52.58 73.33 52.86 ;
      RECT 73.17 52.18 73.33 52.86 ;
      RECT 72.57 51.64 72.73 52.86 ;
      RECT 72.87 12.53 73.03 13.61 ;
      RECT 73.03 11.88 73.19 12.69 ;
      RECT 72.07 11.77 72.31 12.05 ;
      RECT 72.07 11.88 73.19 12.04 ;
      RECT 72.95 8.88 73.11 12.04 ;
      RECT 72.89 62.9 73.05 67.89 ;
      RECT 72.89 65.82 73.11 66.55 ;
      RECT 72.57 47.39 72.73 49.72 ;
      RECT 72.57 47.39 73.05 47.55 ;
      RECT 72.89 43.85 73.05 47.55 ;
      RECT 72.27 43.85 73.05 44.01 ;
      RECT 72.27 39.56 72.43 44.01 ;
      RECT 72.27 39.56 72.61 39.84 ;
      RECT 72.45 39.16 72.61 39.84 ;
      RECT 72.87 22.01 73.03 23.37 ;
      RECT 72.25 22.01 73.03 22.17 ;
      RECT 72.55 24.72 72.93 24.96 ;
      RECT 72.55 22.35 72.71 24.96 ;
      RECT 72.59 34.44 72.93 34.72 ;
      RECT 72.77 32.44 72.93 34.72 ;
      RECT 72.59 33.11 72.93 33.39 ;
      RECT 72.59 32.44 72.93 32.72 ;
      RECT 72.59 40.7 72.93 40.98 ;
      RECT 72.77 38.7 72.93 40.98 ;
      RECT 72.59 40.03 72.93 40.31 ;
      RECT 72.59 38.7 72.93 38.98 ;
      RECT 71.29 12.21 71.45 13.28 ;
      RECT 71.29 12.21 72.87 12.37 ;
      RECT 71.75 11.47 71.91 12.37 ;
      RECT 71.81 10.85 71.97 11.63 ;
      RECT 72.41 62.9 72.57 67.89 ;
      RECT 72.41 64.59 72.69 65.31 ;
      RECT 71.93 46.75 72.09 47.43 ;
      RECT 71.61 46.75 72.41 46.91 ;
      RECT 72.25 44.23 72.41 46.91 ;
      RECT 71.61 44.23 71.77 46.91 ;
      RECT 72.13 10.51 72.29 11.24 ;
      RECT 71.63 10.51 72.29 10.67 ;
      RECT 71.98 8.96 72.14 9.79 ;
      RECT 70.95 8.96 72.14 9.12 ;
      RECT 71.65 20.63 71.93 20.79 ;
      RECT 71.77 19.59 71.93 20.79 ;
      RECT 69.71 34.88 71.91 35.04 ;
      RECT 71.63 34.59 71.91 35.04 ;
      RECT 70.69 34.59 70.93 35.04 ;
      RECT 69.71 34.59 69.99 35.04 ;
      RECT 70.69 38.38 70.93 39.02 ;
      RECT 71.63 38.38 71.91 38.83 ;
      RECT 69.71 38.38 69.99 38.83 ;
      RECT 69.71 38.38 71.91 38.54 ;
      RECT 71.53 28.04 71.85 28.32 ;
      RECT 71.53 25.99 71.69 28.32 ;
      RECT 70.34 27.02 70.5 27.7 ;
      RECT 70.34 27.02 71.69 27.18 ;
      RECT 71.31 25.99 71.69 26.23 ;
      RECT 71.31 25.16 71.47 26.23 ;
      RECT 69.87 36.47 71.75 36.63 ;
      RECT 71.59 35.88 71.75 36.63 ;
      RECT 70.73 35.23 70.89 36.63 ;
      RECT 69.87 35.88 70.03 36.63 ;
      RECT 71.69 35.23 71.85 36.06 ;
      RECT 69.77 35.23 69.93 36.06 ;
      RECT 71.69 37.11 71.85 38.19 ;
      RECT 70.73 36.79 70.89 38.19 ;
      RECT 69.77 37.11 69.93 38.19 ;
      RECT 71.59 36.79 71.75 37.39 ;
      RECT 69.87 36.79 70.03 37.39 ;
      RECT 69.87 36.79 71.75 36.95 ;
      RECT 70.99 22.01 71.15 23.37 ;
      RECT 70.99 22.01 71.77 22.17 ;
      RECT 69.95 68.07 71.77 68.23 ;
      RECT 69.95 62.02 70.11 68.23 ;
      RECT 69.95 62.02 70.33 62.18 ;
      RECT 70.17 57.45 70.33 62.18 ;
      RECT 70.17 57.45 71.77 57.61 ;
      RECT 71.45 57.39 71.77 57.61 ;
      RECT 71.45 53.74 71.61 57.61 ;
      RECT 71.61 51.32 71.77 53.9 ;
      RECT 71.29 51.32 71.77 51.48 ;
      RECT 71.29 49.88 71.45 51.48 ;
      RECT 70.97 49.88 71.45 50.04 ;
      RECT 70.97 47.71 71.13 50.04 ;
      RECT 70.51 47.71 71.13 47.99 ;
      RECT 71.29 47.39 71.45 49.72 ;
      RECT 70.97 47.39 71.45 47.55 ;
      RECT 70.97 43.85 71.13 47.55 ;
      RECT 70.97 43.85 71.75 44.01 ;
      RECT 71.59 39.56 71.75 44.01 ;
      RECT 71.41 39.56 71.75 39.84 ;
      RECT 71.41 39.16 71.57 39.84 ;
      RECT 71.11 14.44 71.27 15.64 ;
      RECT 71.11 14.44 71.61 14.6 ;
      RECT 71.45 62.9 71.61 67.89 ;
      RECT 71.33 64.59 71.61 65.31 ;
      RECT 71.09 24.72 71.47 24.96 ;
      RECT 71.31 22.35 71.47 24.96 ;
      RECT 70.81 12.32 70.97 13.37 ;
      RECT 70.93 11.56 71.09 12.48 ;
      RECT 70.33 11.56 71.45 11.72 ;
      RECT 71.29 10.27 71.45 11.72 ;
      RECT 70.33 10.4 70.49 11.72 ;
      RECT 70.69 52.58 71.45 52.86 ;
      RECT 71.29 51.64 71.45 52.86 ;
      RECT 70.69 52.18 70.85 52.86 ;
      RECT 71.09 34.44 71.43 34.72 ;
      RECT 71.09 32.44 71.25 34.72 ;
      RECT 71.09 33.11 71.43 33.39 ;
      RECT 71.09 32.44 71.43 32.72 ;
      RECT 71.09 40.7 71.43 40.98 ;
      RECT 71.09 38.7 71.25 40.98 ;
      RECT 71.09 40.03 71.43 40.31 ;
      RECT 71.09 38.7 71.43 38.98 ;
      RECT 71.15 53.23 71.43 53.51 ;
      RECT 71.15 53.03 71.31 53.51 ;
      RECT 70.33 53.03 71.31 53.19 ;
      RECT 70.33 50.98 70.49 53.19 ;
      RECT 70.29 52.54 70.49 52.82 ;
      RECT 69.95 50.98 70.49 51.14 ;
      RECT 69.95 50.8 70.17 51.14 ;
      RECT 69.85 56.67 70.01 61.86 ;
      RECT 69.85 56.67 71.29 56.83 ;
      RECT 71.13 56 71.29 56.83 ;
      RECT 70.01 54.4 70.17 56.83 ;
      RECT 70.99 26.36 71.15 26.72 ;
      RECT 68.85 26.36 71.15 26.52 ;
      RECT 68.85 26.04 69.01 26.52 ;
      RECT 68.2 26.04 69.01 26.2 ;
      RECT 70.97 50.66 71.13 51.5 ;
      RECT 70.33 50.66 71.13 50.82 ;
      RECT 70.33 50.18 70.49 50.82 ;
      RECT 69.85 50.18 70.49 50.5 ;
      RECT 69.85 47.07 70.01 50.5 ;
      RECT 69.85 47.07 70.33 47.23 ;
      RECT 70.17 45.44 70.33 47.23 ;
      RECT 70.73 55.68 70.89 56.51 ;
      RECT 70.73 55.68 71.13 55.84 ;
      RECT 70.97 53.67 71.13 55.84 ;
      RECT 70.49 53.67 71.13 53.83 ;
      RECT 70.49 53.35 70.77 53.83 ;
      RECT 70.97 62.9 71.13 67.89 ;
      RECT 70.91 65.82 71.13 66.55 ;
      RECT 70.65 51.7 71.03 51.92 ;
      RECT 70.65 50.98 70.81 51.92 ;
      RECT 68.82 28.01 70.98 28.17 ;
      RECT 70.82 27.34 70.98 28.17 ;
      RECT 70.66 27.93 70.98 28.17 ;
      RECT 69.82 26.97 69.98 28.17 ;
      RECT 68.82 26.68 68.98 28.17 ;
      RECT 70.33 12 70.49 12.84 ;
      RECT 70.33 12 70.77 12.16 ;
      RECT 70.61 11.88 70.77 12.16 ;
      RECT 69.08 8.82 70.67 8.98 ;
      RECT 70.51 7.16 70.67 8.98 ;
      RECT 70.17 47.39 70.33 49.72 ;
      RECT 70.17 47.39 70.65 47.55 ;
      RECT 70.49 43.85 70.65 47.55 ;
      RECT 69.87 43.85 70.65 44.01 ;
      RECT 69.87 39.56 70.03 44.01 ;
      RECT 69.87 39.56 70.21 39.84 ;
      RECT 70.05 39.16 70.21 39.84 ;
      RECT 70.48 9.92 70.64 10.24 ;
      RECT 70.24 9.92 70.64 10.12 ;
      RECT 69.45 15.8 69.61 17.77 ;
      RECT 69.45 15.8 70.27 15.96 ;
      RECT 70.27 14.42 70.43 15.88 ;
      RECT 70.09 15.72 70.43 15.88 ;
      RECT 70.27 14.42 70.61 14.58 ;
      RECT 70.33 24.79 70.53 25.35 ;
      RECT 70.21 24.79 70.53 25.03 ;
      RECT 70.19 34.44 70.53 34.72 ;
      RECT 70.37 32.44 70.53 34.72 ;
      RECT 70.19 33.11 70.53 33.39 ;
      RECT 70.19 32.44 70.53 32.72 ;
      RECT 70.19 40.7 70.53 40.98 ;
      RECT 70.37 38.7 70.53 40.98 ;
      RECT 70.19 40.03 70.53 40.31 ;
      RECT 70.19 38.7 70.53 38.98 ;
      RECT 70.21 21.85 70.37 24.3 ;
      RECT 70.21 21.85 70.51 22.13 ;
      RECT 70.33 54.06 70.49 56.51 ;
      RECT 69.97 54.06 70.49 54.22 ;
      RECT 69.97 52.98 70.17 54.22 ;
      RECT 69.97 51.34 70.13 54.22 ;
      RECT 69.97 51.34 70.17 52.12 ;
      RECT 69.83 18.51 70.02 18.94 ;
      RECT 69.63 18.51 70.32 18.7 ;
      RECT 69.81 21.29 69.97 23.37 ;
      RECT 69.89 19.81 70.05 21.46 ;
      RECT 69.43 12.58 69.71 13.24 ;
      RECT 69.55 11.84 69.71 13.24 ;
      RECT 69.19 11.84 69.35 12.12 ;
      RECT 69.19 11.84 70.03 12 ;
      RECT 69.87 10.46 70.03 12 ;
      RECT 69.53 46.75 69.69 47.43 ;
      RECT 69.21 46.75 70.01 46.91 ;
      RECT 69.85 44.23 70.01 46.91 ;
      RECT 69.21 44.23 69.37 46.91 ;
      RECT 69.37 26.02 69.93 26.18 ;
      RECT 69.37 25.58 69.53 26.18 ;
      RECT 68.83 25.58 69.53 25.74 ;
      RECT 68.83 24 69.03 25.74 ;
      RECT 68.09 24.24 69.03 24.52 ;
      RECT 68.09 21.85 68.25 24.52 ;
      RECT 68.76 9.14 68.95 9.52 ;
      RECT 68.76 9.14 69.89 9.3 ;
      RECT 68.76 8.52 68.92 9.52 ;
      RECT 68.74 8.36 68.9 8.64 ;
      RECT 69.13 18.13 69.79 18.3 ;
      RECT 69.13 15 69.29 18.3 ;
      RECT 69.13 15.32 69.83 15.64 ;
      RECT 68.67 15 69.29 15.16 ;
      RECT 69.39 9.68 69.55 11.68 ;
      RECT 64.87 9.68 65.03 11.68 ;
      RECT 67.93 9.68 68.09 11.36 ;
      RECT 66.33 9.68 66.49 11.36 ;
      RECT 66.33 10.76 68.09 10.92 ;
      RECT 67.13 8.38 67.29 10.92 ;
      RECT 67.93 9.68 69.55 9.84 ;
      RECT 69.27 9.46 69.43 9.84 ;
      RECT 64.87 9.68 66.49 9.84 ;
      RECT 64.99 9.46 65.15 9.84 ;
      RECT 69.34 26.68 69.5 27.85 ;
      RECT 69.3 26.68 69.54 27.33 ;
      RECT 67.31 34.88 69.51 35.04 ;
      RECT 69.23 34.59 69.51 35.04 ;
      RECT 68.29 34.59 68.53 35.04 ;
      RECT 67.31 34.59 67.59 35.04 ;
      RECT 68.29 38.38 68.53 39.02 ;
      RECT 69.23 38.38 69.51 38.83 ;
      RECT 67.31 38.38 67.59 38.83 ;
      RECT 67.31 38.38 69.51 38.54 ;
      RECT 69.29 13.5 69.45 14.2 ;
      RECT 69.11 13.5 69.45 13.66 ;
      RECT 69.11 12.52 69.27 13.66 ;
      RECT 68.87 12.52 69.27 12.84 ;
      RECT 68.87 10.84 69.03 12.84 ;
      RECT 67.47 36.47 69.35 36.63 ;
      RECT 69.19 35.86 69.35 36.63 ;
      RECT 68.33 35.23 68.49 36.63 ;
      RECT 67.47 35.86 67.63 36.63 ;
      RECT 69.29 35.23 69.45 36.05 ;
      RECT 67.37 35.23 67.53 36.05 ;
      RECT 69.29 37.11 69.45 38.19 ;
      RECT 68.33 36.79 68.49 38.19 ;
      RECT 67.37 37.11 67.53 38.19 ;
      RECT 69.19 36.79 69.35 37.39 ;
      RECT 67.47 36.79 67.63 37.39 ;
      RECT 67.47 36.79 69.35 36.95 ;
      RECT 68.09 50.66 68.25 51.5 ;
      RECT 68.09 50.66 68.89 50.82 ;
      RECT 68.73 50.18 68.89 50.82 ;
      RECT 68.73 50.18 69.37 50.5 ;
      RECT 69.21 47.07 69.37 50.5 ;
      RECT 68.89 47.07 69.37 47.23 ;
      RECT 68.89 45.44 69.05 47.23 ;
      RECT 69.21 56.67 69.37 61.86 ;
      RECT 67.93 56.67 69.37 56.83 ;
      RECT 69.05 54.4 69.21 56.83 ;
      RECT 67.93 56 68.09 56.83 ;
      RECT 68.89 47.39 69.05 49.72 ;
      RECT 68.57 47.39 69.05 47.55 ;
      RECT 68.57 43.85 68.73 47.55 ;
      RECT 68.57 43.85 69.35 44.01 ;
      RECT 69.19 39.56 69.35 44.01 ;
      RECT 69.01 39.56 69.35 39.84 ;
      RECT 69.01 39.16 69.17 39.84 ;
      RECT 69.15 23.12 69.31 23.84 ;
      RECT 68.41 23.12 69.31 23.28 ;
      RECT 68.41 20.86 68.57 23.28 ;
      RECT 68.41 20.86 68.77 21.02 ;
      RECT 68.61 20.74 68.77 21.02 ;
      RECT 67.8 28.52 68.89 28.68 ;
      RECT 68.61 28.35 68.89 28.68 ;
      RECT 68.61 28.35 69.29 28.51 ;
      RECT 67.79 53.23 68.07 53.51 ;
      RECT 67.91 53.03 68.07 53.51 ;
      RECT 67.91 53.03 68.89 53.19 ;
      RECT 68.73 50.98 68.89 53.19 ;
      RECT 68.73 52.54 68.93 52.82 ;
      RECT 68.73 50.98 69.27 51.14 ;
      RECT 69.05 50.8 69.27 51.14 ;
      RECT 67.45 68.07 69.27 68.23 ;
      RECT 69.11 62.02 69.27 68.23 ;
      RECT 68.89 62.02 69.27 62.18 ;
      RECT 68.89 57.45 69.05 62.18 ;
      RECT 67.45 57.45 69.05 57.61 ;
      RECT 67.45 57.39 67.77 57.61 ;
      RECT 67.61 53.74 67.77 57.61 ;
      RECT 67.45 51.32 67.61 53.9 ;
      RECT 67.45 51.32 67.93 51.48 ;
      RECT 67.77 49.88 67.93 51.48 ;
      RECT 67.77 49.88 68.25 50.04 ;
      RECT 68.09 47.71 68.25 50.04 ;
      RECT 68.09 47.71 68.71 47.99 ;
      RECT 68.73 54.06 68.89 56.51 ;
      RECT 68.73 54.06 69.25 54.22 ;
      RECT 69.09 51.34 69.25 54.22 ;
      RECT 69.05 52.98 69.25 54.22 ;
      RECT 69.05 51.34 69.25 52.12 ;
      RECT 68.69 13.06 68.85 13.54 ;
      RECT 68.41 13.06 68.85 13.22 ;
      RECT 68.41 10 68.57 13.22 ;
      RECT 68.41 10 69.23 10.16 ;
      RECT 68.77 22.29 69.01 22.53 ;
      RECT 68.77 21.18 68.93 22.53 ;
      RECT 68.73 21.18 68.93 21.58 ;
      RECT 68.93 19.81 69.1 21.35 ;
      RECT 68.69 34.44 69.03 34.72 ;
      RECT 68.69 32.44 68.85 34.72 ;
      RECT 68.69 33.11 69.03 33.39 ;
      RECT 68.69 32.44 69.03 32.72 ;
      RECT 68.69 40.7 69.03 40.98 ;
      RECT 68.69 38.7 68.85 40.98 ;
      RECT 68.69 40.03 69.03 40.31 ;
      RECT 68.69 38.7 69.03 38.98 ;
      RECT 68.57 17.24 68.73 19 ;
      RECT 67.61 14.39 67.77 18.85 ;
      RECT 67.61 17.24 68.73 17.4 ;
      RECT 67.59 15.32 67.79 16.04 ;
      RECT 67.61 14.39 67.79 16.04 ;
      RECT 68.33 55.68 68.49 56.51 ;
      RECT 68.09 55.68 68.49 55.84 ;
      RECT 68.09 53.67 68.25 55.84 ;
      RECT 68.09 53.67 68.73 53.83 ;
      RECT 68.45 53.35 68.73 53.83 ;
      RECT 67.88 24.7 68.04 28.32 ;
      RECT 67.88 25.16 68.57 25.32 ;
      RECT 67.35 24.7 68.04 24.86 ;
      RECT 68.19 51.7 68.57 51.92 ;
      RECT 68.41 50.98 68.57 51.92 ;
      RECT 67.77 52.58 68.53 52.86 ;
      RECT 68.37 52.18 68.53 52.86 ;
      RECT 67.77 51.64 67.93 52.86 ;
      RECT 68.09 62.9 68.25 67.89 ;
      RECT 68.09 65.82 68.31 66.55 ;
      RECT 67.53 9.36 67.69 10.6 ;
      RECT 67.53 9.36 68.27 9.52 ;
      RECT 67.77 47.39 67.93 49.72 ;
      RECT 67.77 47.39 68.25 47.55 ;
      RECT 68.09 43.85 68.25 47.55 ;
      RECT 67.47 43.85 68.25 44.01 ;
      RECT 67.47 39.56 67.63 44.01 ;
      RECT 67.47 39.56 67.81 39.84 ;
      RECT 67.65 39.16 67.81 39.84 ;
      RECT 67.79 34.44 68.13 34.72 ;
      RECT 67.97 32.44 68.13 34.72 ;
      RECT 67.79 33.11 68.13 33.39 ;
      RECT 67.79 32.44 68.13 32.72 ;
      RECT 67.79 40.7 68.13 40.98 ;
      RECT 67.97 38.7 68.13 40.98 ;
      RECT 67.79 40.03 68.13 40.31 ;
      RECT 67.79 38.7 68.13 38.98 ;
      RECT 67.69 11.52 67.85 12.43 ;
      RECT 67.69 11.75 67.93 12.03 ;
      RECT 67.41 11.52 67.85 11.68 ;
      RECT 67.41 11.08 67.57 11.68 ;
      RECT 67.61 62.9 67.77 67.89 ;
      RECT 67.61 64.59 67.89 65.31 ;
      RECT 67.61 23.73 67.79 24.54 ;
      RECT 67.61 20.48 67.77 24.54 ;
      RECT 67.13 46.75 67.29 47.43 ;
      RECT 66.81 46.75 67.61 46.91 ;
      RECT 67.45 44.23 67.61 46.91 ;
      RECT 66.81 44.23 66.97 46.91 ;
      RECT 67.4 26.15 67.56 28.96 ;
      RECT 67.37 26.15 67.56 26.51 ;
      RECT 64.91 34.88 67.11 35.04 ;
      RECT 66.83 34.59 67.11 35.04 ;
      RECT 65.89 34.59 66.13 35.04 ;
      RECT 64.91 34.59 65.19 35.04 ;
      RECT 65.89 38.38 66.13 39.02 ;
      RECT 66.83 38.38 67.11 38.83 ;
      RECT 64.91 38.38 65.19 38.83 ;
      RECT 64.91 38.38 67.11 38.54 ;
      RECT 66.38 24.7 66.54 28.32 ;
      RECT 65.85 25.16 66.54 25.32 ;
      RECT 66.38 24.7 67.07 24.86 ;
      RECT 66.86 26.15 67.02 28.96 ;
      RECT 66.86 26.15 67.05 26.51 ;
      RECT 65.07 36.47 66.95 36.63 ;
      RECT 66.79 35.88 66.95 36.63 ;
      RECT 65.93 35.23 66.09 36.63 ;
      RECT 65.07 35.88 65.23 36.63 ;
      RECT 66.89 35.23 67.05 36.06 ;
      RECT 64.97 35.23 65.13 36.06 ;
      RECT 66.89 37.11 67.05 38.19 ;
      RECT 65.93 36.79 66.09 38.19 ;
      RECT 64.97 37.11 65.13 38.19 ;
      RECT 66.79 36.79 66.95 37.39 ;
      RECT 65.07 36.79 65.23 37.39 ;
      RECT 65.07 36.79 66.95 36.95 ;
      RECT 66.57 11.52 66.73 12.43 ;
      RECT 66.49 11.75 66.73 12.03 ;
      RECT 66.57 11.52 67.01 11.68 ;
      RECT 66.85 11.08 67.01 11.68 ;
      RECT 65.15 68.07 66.97 68.23 ;
      RECT 65.15 62.02 65.31 68.23 ;
      RECT 65.15 62.02 65.53 62.18 ;
      RECT 65.37 57.45 65.53 62.18 ;
      RECT 65.37 57.45 66.97 57.61 ;
      RECT 66.65 57.39 66.97 57.61 ;
      RECT 66.65 53.74 66.81 57.61 ;
      RECT 66.81 51.32 66.97 53.9 ;
      RECT 66.49 51.32 66.97 51.48 ;
      RECT 66.49 49.88 66.65 51.48 ;
      RECT 66.17 49.88 66.65 50.04 ;
      RECT 66.17 47.71 66.33 50.04 ;
      RECT 65.71 47.71 66.33 47.99 ;
      RECT 66.49 47.39 66.65 49.72 ;
      RECT 66.17 47.39 66.65 47.55 ;
      RECT 66.17 43.85 66.33 47.55 ;
      RECT 66.17 43.85 66.95 44.01 ;
      RECT 66.79 39.56 66.95 44.01 ;
      RECT 66.61 39.56 66.95 39.84 ;
      RECT 66.61 39.16 66.77 39.84 ;
      RECT 66.73 9.36 66.89 10.6 ;
      RECT 66.15 9.36 66.89 9.52 ;
      RECT 65.69 17.24 65.85 19 ;
      RECT 66.65 14.39 66.81 18.85 ;
      RECT 65.69 17.24 66.81 17.4 ;
      RECT 66.63 15.32 66.83 16.04 ;
      RECT 66.63 14.39 66.81 16.04 ;
      RECT 66.63 23.73 66.81 24.54 ;
      RECT 66.65 20.48 66.81 24.54 ;
      RECT 66.65 62.9 66.81 67.89 ;
      RECT 66.53 64.59 66.81 65.31 ;
      RECT 65.89 52.58 66.65 52.86 ;
      RECT 66.49 51.64 66.65 52.86 ;
      RECT 65.89 52.18 66.05 52.86 ;
      RECT 66.29 34.44 66.63 34.72 ;
      RECT 66.29 32.44 66.45 34.72 ;
      RECT 66.29 33.11 66.63 33.39 ;
      RECT 66.29 32.44 66.63 32.72 ;
      RECT 66.29 40.7 66.63 40.98 ;
      RECT 66.29 38.7 66.45 40.98 ;
      RECT 66.29 40.03 66.63 40.31 ;
      RECT 66.29 38.7 66.63 38.98 ;
      RECT 66.35 53.23 66.63 53.51 ;
      RECT 66.35 53.03 66.51 53.51 ;
      RECT 65.53 53.03 66.51 53.19 ;
      RECT 65.53 50.98 65.69 53.19 ;
      RECT 65.49 52.54 65.69 52.82 ;
      RECT 65.15 50.98 65.69 51.14 ;
      RECT 65.15 50.8 65.37 51.14 ;
      RECT 65.53 28.52 66.62 28.68 ;
      RECT 65.53 28.35 65.81 28.68 ;
      RECT 65.13 28.35 65.81 28.51 ;
      RECT 65.05 56.67 65.21 61.86 ;
      RECT 65.05 56.67 66.49 56.83 ;
      RECT 66.33 56 66.49 56.83 ;
      RECT 65.21 54.4 65.37 56.83 ;
      RECT 64.49 26.02 65.05 26.18 ;
      RECT 64.89 25.58 65.05 26.18 ;
      RECT 64.89 25.58 65.59 25.74 ;
      RECT 65.39 24 65.59 25.74 ;
      RECT 65.39 24.24 66.33 24.52 ;
      RECT 66.17 21.85 66.33 24.52 ;
      RECT 66.17 50.66 66.33 51.5 ;
      RECT 65.53 50.66 66.33 50.82 ;
      RECT 65.53 50.18 65.69 50.82 ;
      RECT 65.05 50.18 65.69 50.5 ;
      RECT 65.05 47.07 65.21 50.5 ;
      RECT 65.05 47.07 65.53 47.23 ;
      RECT 65.37 45.44 65.53 47.23 ;
      RECT 65.93 55.68 66.09 56.51 ;
      RECT 65.93 55.68 66.33 55.84 ;
      RECT 66.17 53.67 66.33 55.84 ;
      RECT 65.69 53.67 66.33 53.83 ;
      RECT 65.69 53.35 65.97 53.83 ;
      RECT 66.17 62.9 66.33 67.89 ;
      RECT 66.11 65.82 66.33 66.55 ;
      RECT 65.85 51.7 66.23 51.92 ;
      RECT 65.85 50.98 66.01 51.92 ;
      RECT 63.27 26.36 63.43 26.72 ;
      RECT 63.27 26.36 65.57 26.52 ;
      RECT 65.41 26.04 65.57 26.52 ;
      RECT 65.41 26.04 66.22 26.2 ;
      RECT 65.57 13.06 65.73 13.54 ;
      RECT 65.57 13.06 66.01 13.22 ;
      RECT 65.85 10 66.01 13.22 ;
      RECT 65.19 10 66.01 10.16 ;
      RECT 65.11 23.12 65.27 23.84 ;
      RECT 65.11 23.12 66.01 23.28 ;
      RECT 65.85 20.86 66.01 23.28 ;
      RECT 65.65 20.86 66.01 21.02 ;
      RECT 65.65 20.74 65.81 21.02 ;
      RECT 65.37 47.39 65.53 49.72 ;
      RECT 65.37 47.39 65.85 47.55 ;
      RECT 65.69 43.85 65.85 47.55 ;
      RECT 65.07 43.85 65.85 44.01 ;
      RECT 65.07 39.56 65.23 44.01 ;
      RECT 65.07 39.56 65.41 39.84 ;
      RECT 65.25 39.16 65.41 39.84 ;
      RECT 64.63 18.13 65.29 18.3 ;
      RECT 65.13 15 65.29 18.3 ;
      RECT 64.59 15.32 65.29 15.64 ;
      RECT 65.13 15 65.75 15.16 ;
      RECT 65.39 34.44 65.73 34.72 ;
      RECT 65.57 32.44 65.73 34.72 ;
      RECT 65.39 33.11 65.73 33.39 ;
      RECT 65.39 32.44 65.73 32.72 ;
      RECT 65.39 40.7 65.73 40.98 ;
      RECT 65.57 38.7 65.73 40.98 ;
      RECT 65.39 40.03 65.73 40.31 ;
      RECT 65.39 38.7 65.73 38.98 ;
      RECT 65.41 22.29 65.65 22.53 ;
      RECT 65.49 21.18 65.65 22.53 ;
      RECT 65.49 21.18 65.69 21.58 ;
      RECT 65.32 19.81 65.49 21.35 ;
      RECT 65.53 54.06 65.69 56.51 ;
      RECT 65.17 54.06 65.69 54.22 ;
      RECT 65.17 52.98 65.37 54.22 ;
      RECT 65.17 51.34 65.33 54.22 ;
      RECT 65.17 51.34 65.37 52.12 ;
      RECT 65.47 9.14 65.66 9.52 ;
      RECT 64.53 9.14 65.66 9.3 ;
      RECT 65.5 8.52 65.66 9.52 ;
      RECT 65.52 8.36 65.68 8.64 ;
      RECT 63.44 28.01 65.6 28.17 ;
      RECT 65.44 26.68 65.6 28.17 ;
      RECT 64.44 26.97 64.6 28.17 ;
      RECT 63.44 27.93 63.76 28.17 ;
      RECT 63.44 27.34 63.6 28.17 ;
      RECT 64.97 13.5 65.13 14.2 ;
      RECT 64.97 13.5 65.31 13.66 ;
      RECT 65.15 12.52 65.31 13.66 ;
      RECT 65.15 12.52 65.55 12.84 ;
      RECT 65.39 10.84 65.55 12.84 ;
      RECT 63.75 8.82 65.34 8.98 ;
      RECT 63.75 7.16 63.91 8.98 ;
      RECT 64.71 12.58 64.99 13.24 ;
      RECT 64.71 11.84 64.87 13.24 ;
      RECT 65.07 11.84 65.23 12.12 ;
      RECT 64.39 11.84 65.23 12 ;
      RECT 64.39 10.46 64.55 12 ;
      RECT 64.73 46.75 64.89 47.43 ;
      RECT 64.41 46.75 65.21 46.91 ;
      RECT 65.05 44.23 65.21 46.91 ;
      RECT 64.41 44.23 64.57 46.91 ;
      RECT 64.92 26.68 65.08 27.85 ;
      RECT 64.88 26.68 65.12 27.33 ;
      RECT 64.81 15.8 64.97 17.77 ;
      RECT 64.15 15.8 64.97 15.96 ;
      RECT 63.99 14.42 64.15 15.88 ;
      RECT 63.99 15.72 64.33 15.88 ;
      RECT 63.81 14.42 64.15 14.58 ;
      RECT 59.85 28.74 64.97 28.9 ;
      RECT 63.05 27.92 63.21 28.9 ;
      RECT 61.61 27.92 61.77 28.9 ;
      RECT 64.4 18.51 64.59 18.94 ;
      RECT 64.1 18.51 64.79 18.7 ;
      RECT 62.51 34.88 64.71 35.04 ;
      RECT 64.43 34.59 64.71 35.04 ;
      RECT 63.49 34.59 63.73 35.04 ;
      RECT 62.51 34.59 62.79 35.04 ;
      RECT 63.49 38.38 63.73 39.02 ;
      RECT 64.43 38.38 64.71 38.83 ;
      RECT 62.51 38.38 62.79 38.83 ;
      RECT 62.51 38.38 64.71 38.54 ;
      RECT 62.33 21.69 62.49 26.21 ;
      RECT 63.57 24.35 63.73 26.2 ;
      RECT 61.09 24.34 61.25 26.2 ;
      RECT 64.45 24.04 64.67 25.52 ;
      RECT 60.15 24.04 60.37 25.52 ;
      RECT 63.57 24.46 64.67 24.63 ;
      RECT 60.15 24.46 61.25 24.63 ;
      RECT 61.07 21.69 61.23 24.63 ;
      RECT 63.59 21.69 63.75 24.63 ;
      RECT 61.07 21.69 63.75 21.85 ;
      RECT 60.56 18.78 61.68 18.94 ;
      RECT 63.44 16.44 63.6 18.8 ;
      RECT 62.47 17.26 62.64 18.8 ;
      RECT 61.52 16.03 61.68 18.94 ;
      RECT 60.56 17.48 60.74 18.94 ;
      RECT 63.44 16.44 63.65 17.57 ;
      RECT 60.58 16.44 60.74 18.94 ;
      RECT 62.47 17.26 63.65 17.42 ;
      RECT 63.37 16.44 63.65 17.42 ;
      RECT 62.47 16.12 62.63 18.8 ;
      RECT 60.71 14.52 60.87 16.71 ;
      RECT 61.52 16.12 64.65 16.28 ;
      RECT 62.67 14.84 62.83 16.28 ;
      RECT 61.67 14.52 61.83 16.28 ;
      RECT 60.71 14.52 61.83 14.68 ;
      RECT 62.67 36.47 64.55 36.63 ;
      RECT 64.39 35.86 64.55 36.63 ;
      RECT 63.53 35.23 63.69 36.63 ;
      RECT 62.67 35.86 62.83 36.63 ;
      RECT 64.49 35.23 64.65 36.05 ;
      RECT 62.57 35.23 62.73 36.05 ;
      RECT 64.49 37.11 64.65 38.19 ;
      RECT 63.53 36.79 63.69 38.19 ;
      RECT 62.57 37.11 62.73 38.19 ;
      RECT 64.39 36.79 64.55 37.39 ;
      RECT 62.67 36.79 62.83 37.39 ;
      RECT 62.67 36.79 64.55 36.95 ;
      RECT 64.45 21.29 64.61 23.37 ;
      RECT 64.37 19.81 64.53 21.46 ;
      RECT 63.29 50.66 63.45 51.5 ;
      RECT 63.29 50.66 64.09 50.82 ;
      RECT 63.93 50.18 64.09 50.82 ;
      RECT 63.93 50.18 64.57 50.5 ;
      RECT 64.41 47.07 64.57 50.5 ;
      RECT 64.09 47.07 64.57 47.23 ;
      RECT 64.09 45.44 64.25 47.23 ;
      RECT 64.41 56.67 64.57 61.86 ;
      RECT 63.13 56.67 64.57 56.83 ;
      RECT 64.25 54.4 64.41 56.83 ;
      RECT 63.13 56 63.29 56.83 ;
      RECT 64.09 47.39 64.25 49.72 ;
      RECT 63.77 47.39 64.25 47.55 ;
      RECT 63.77 43.85 63.93 47.55 ;
      RECT 63.77 43.85 64.55 44.01 ;
      RECT 64.39 39.56 64.55 44.01 ;
      RECT 64.21 39.56 64.55 39.84 ;
      RECT 64.21 39.16 64.37 39.84 ;
      RECT 62.99 53.23 63.27 53.51 ;
      RECT 63.11 53.03 63.27 53.51 ;
      RECT 63.11 53.03 64.09 53.19 ;
      RECT 63.93 50.98 64.09 53.19 ;
      RECT 63.93 52.54 64.13 52.82 ;
      RECT 63.93 50.98 64.47 51.14 ;
      RECT 64.25 50.8 64.47 51.14 ;
      RECT 62.65 68.07 64.47 68.23 ;
      RECT 64.31 62.02 64.47 68.23 ;
      RECT 64.09 62.02 64.47 62.18 ;
      RECT 64.09 57.45 64.25 62.18 ;
      RECT 62.65 57.45 64.25 57.61 ;
      RECT 62.65 57.39 62.97 57.61 ;
      RECT 62.81 53.74 62.97 57.61 ;
      RECT 62.65 51.32 62.81 53.9 ;
      RECT 62.65 51.32 63.13 51.48 ;
      RECT 62.97 49.88 63.13 51.48 ;
      RECT 62.97 49.88 63.45 50.04 ;
      RECT 63.29 47.71 63.45 50.04 ;
      RECT 63.29 47.71 63.91 47.99 ;
      RECT 63.93 54.06 64.09 56.51 ;
      RECT 63.93 54.06 64.45 54.22 ;
      RECT 64.29 51.34 64.45 54.22 ;
      RECT 64.25 52.98 64.45 54.22 ;
      RECT 64.25 51.34 64.45 52.12 ;
      RECT 63.89 34.44 64.23 34.72 ;
      RECT 63.89 32.44 64.05 34.72 ;
      RECT 63.89 33.11 64.23 33.39 ;
      RECT 63.89 32.44 64.23 32.72 ;
      RECT 63.89 40.7 64.23 40.98 ;
      RECT 63.89 38.7 64.05 40.98 ;
      RECT 63.89 40.03 64.23 40.31 ;
      RECT 63.89 38.7 64.23 38.98 ;
      RECT 60.21 21.37 60.37 23.37 ;
      RECT 60.21 21.37 64.21 21.53 ;
      RECT 64.05 20.78 64.21 21.53 ;
      RECT 60.7 20.73 60.86 21.53 ;
      RECT 64.05 21.85 64.21 24.3 ;
      RECT 63.91 21.85 64.21 22.13 ;
      RECT 63.89 24.79 64.09 25.35 ;
      RECT 63.89 24.79 64.21 25.03 ;
      RECT 63.78 9.92 63.94 10.24 ;
      RECT 63.78 9.92 64.18 10.12 ;
      RECT 63.45 12.32 63.61 13.37 ;
      RECT 63.33 11.56 63.49 12.48 ;
      RECT 62.97 11.56 64.09 11.72 ;
      RECT 63.93 10.4 64.09 11.72 ;
      RECT 62.97 10.27 63.13 11.72 ;
      RECT 63.93 12 64.09 12.84 ;
      RECT 63.65 12 64.09 12.16 ;
      RECT 63.65 11.88 63.81 12.16 ;
      RECT 62.57 28.04 62.89 28.32 ;
      RECT 62.73 25.99 62.89 28.32 ;
      RECT 63.92 27.02 64.08 27.7 ;
      RECT 62.73 27.02 64.08 27.18 ;
      RECT 62.73 25.99 63.11 26.23 ;
      RECT 62.95 25.16 63.11 26.23 ;
      RECT 63.53 55.68 63.69 56.51 ;
      RECT 63.29 55.68 63.69 55.84 ;
      RECT 63.29 53.67 63.45 55.84 ;
      RECT 63.29 53.67 63.93 53.83 ;
      RECT 63.65 53.35 63.93 53.83 ;
      RECT 63.39 51.7 63.77 51.92 ;
      RECT 63.61 50.98 63.77 51.92 ;
      RECT 62.97 52.58 63.73 52.86 ;
      RECT 63.57 52.18 63.73 52.86 ;
      RECT 62.97 51.64 63.13 52.86 ;
      RECT 61.79 8.5 61.95 11.72 ;
      RECT 60.83 8.12 60.99 11.72 ;
      RECT 59.87 9.28 60.03 11.72 ;
      RECT 63.45 9.63 63.61 11.4 ;
      RECT 61.79 9.95 63.61 10.11 ;
      RECT 62.76 9.79 62.92 10.11 ;
      RECT 59.79 8.12 59.99 9.84 ;
      RECT 63.16 9.63 63.67 9.79 ;
      RECT 59.79 9.28 60.99 9.44 ;
      RECT 61.68 8.5 61.99 8.78 ;
      RECT 60.83 8.56 61.99 8.72 ;
      RECT 63.29 62.9 63.45 67.89 ;
      RECT 63.29 65.82 63.51 66.55 ;
      RECT 62.28 8.96 62.44 9.79 ;
      RECT 62.28 8.96 63.47 9.12 ;
      RECT 62.97 47.39 63.13 49.72 ;
      RECT 62.97 47.39 63.45 47.55 ;
      RECT 63.29 43.85 63.45 47.55 ;
      RECT 62.67 43.85 63.45 44.01 ;
      RECT 62.67 39.56 62.83 44.01 ;
      RECT 62.67 39.56 63.01 39.84 ;
      RECT 62.85 39.16 63.01 39.84 ;
      RECT 63.27 22.01 63.43 23.37 ;
      RECT 62.65 22.01 63.43 22.17 ;
      RECT 62.95 24.72 63.33 24.96 ;
      RECT 62.95 22.35 63.11 24.96 ;
      RECT 62.99 34.44 63.33 34.72 ;
      RECT 63.17 32.44 63.33 34.72 ;
      RECT 62.99 33.11 63.33 33.39 ;
      RECT 62.99 32.44 63.33 32.72 ;
      RECT 62.99 40.7 63.33 40.98 ;
      RECT 63.17 38.7 63.33 40.98 ;
      RECT 62.99 40.03 63.33 40.31 ;
      RECT 62.99 38.7 63.33 38.98 ;
      RECT 63.15 14.44 63.31 15.64 ;
      RECT 62.81 14.44 63.31 14.6 ;
      RECT 62.97 12.21 63.13 13.28 ;
      RECT 61.55 12.21 63.13 12.37 ;
      RECT 62.51 11.47 62.67 12.37 ;
      RECT 62.45 10.85 62.61 11.63 ;
      RECT 62.81 62.9 62.97 67.89 ;
      RECT 62.81 64.59 63.09 65.31 ;
      RECT 62.33 46.75 62.49 47.43 ;
      RECT 62.01 46.75 62.81 46.91 ;
      RECT 62.65 44.23 62.81 46.91 ;
      RECT 62.01 44.23 62.17 46.91 ;
      RECT 62.13 10.51 62.29 11.24 ;
      RECT 62.13 10.51 62.79 10.67 ;
      RECT 62.49 20.63 62.77 20.79 ;
      RECT 62.49 19.59 62.65 20.79 ;
      RECT 61.39 12.53 61.55 13.61 ;
      RECT 61.23 11.88 61.39 12.69 ;
      RECT 62.11 11.77 62.35 12.05 ;
      RECT 61.23 11.88 62.35 12.04 ;
      RECT 61.31 8.88 61.47 12.04 ;
      RECT 60.11 34.88 62.31 35.04 ;
      RECT 62.03 34.59 62.31 35.04 ;
      RECT 61.09 34.59 61.33 35.04 ;
      RECT 60.11 34.59 60.39 35.04 ;
      RECT 61.09 38.38 61.33 39.02 ;
      RECT 62.03 38.38 62.31 38.83 ;
      RECT 60.11 38.38 60.39 38.83 ;
      RECT 60.11 38.38 62.31 38.54 ;
      RECT 61.93 28.04 62.25 28.32 ;
      RECT 61.93 25.99 62.09 28.32 ;
      RECT 60.74 27.02 60.9 27.7 ;
      RECT 60.74 27.02 62.09 27.18 ;
      RECT 61.71 25.99 62.09 26.23 ;
      RECT 61.71 25.16 61.87 26.23 ;
      RECT 60.27 36.47 62.15 36.63 ;
      RECT 61.99 35.88 62.15 36.63 ;
      RECT 61.13 35.23 61.29 36.63 ;
      RECT 60.27 35.88 60.43 36.63 ;
      RECT 62.09 35.23 62.25 36.06 ;
      RECT 60.17 35.23 60.33 36.06 ;
      RECT 62.09 37.11 62.25 38.19 ;
      RECT 61.13 36.79 61.29 38.19 ;
      RECT 60.17 37.11 60.33 38.19 ;
      RECT 61.99 36.79 62.15 37.39 ;
      RECT 60.27 36.79 60.43 37.39 ;
      RECT 60.27 36.79 62.15 36.95 ;
      RECT 62.07 20.26 62.23 21.05 ;
      RECT 61.5 20.26 62.23 20.44 ;
      RECT 61.5 19.89 61.66 20.44 ;
      RECT 60.84 19.89 61.66 20.05 ;
      RECT 60.84 19.61 61.03 20.05 ;
      RECT 60.75 19.61 61.03 19.77 ;
      RECT 61.39 22.01 61.55 23.37 ;
      RECT 61.39 22.01 62.17 22.17 ;
      RECT 60.35 68.07 62.17 68.23 ;
      RECT 60.35 62.02 60.51 68.23 ;
      RECT 60.35 62.02 60.73 62.18 ;
      RECT 60.57 57.45 60.73 62.18 ;
      RECT 60.57 57.45 62.17 57.61 ;
      RECT 61.85 57.39 62.17 57.61 ;
      RECT 61.85 53.74 62.01 57.61 ;
      RECT 62.01 51.32 62.17 53.9 ;
      RECT 61.69 51.32 62.17 51.48 ;
      RECT 61.69 49.88 61.85 51.48 ;
      RECT 61.37 49.88 61.85 50.04 ;
      RECT 61.37 47.71 61.53 50.04 ;
      RECT 60.91 47.71 61.53 47.99 ;
      RECT 61.69 47.39 61.85 49.72 ;
      RECT 61.37 47.39 61.85 47.55 ;
      RECT 61.37 43.85 61.53 47.55 ;
      RECT 61.37 43.85 62.15 44.01 ;
      RECT 61.99 39.56 62.15 44.01 ;
      RECT 61.81 39.56 62.15 39.84 ;
      RECT 61.81 39.16 61.97 39.84 ;
      RECT 61.85 62.9 62.01 67.89 ;
      RECT 61.73 64.59 62.01 65.31 ;
      RECT 61.49 24.72 61.87 24.96 ;
      RECT 61.71 22.35 61.87 24.96 ;
      RECT 61.09 52.58 61.85 52.86 ;
      RECT 61.69 51.64 61.85 52.86 ;
      RECT 61.09 52.18 61.25 52.86 ;
      RECT 61.49 34.44 61.83 34.72 ;
      RECT 61.49 32.44 61.65 34.72 ;
      RECT 61.49 33.11 61.83 33.39 ;
      RECT 61.49 32.44 61.83 32.72 ;
      RECT 61.49 40.7 61.83 40.98 ;
      RECT 61.49 38.7 61.65 40.98 ;
      RECT 61.49 40.03 61.83 40.31 ;
      RECT 61.49 38.7 61.83 38.98 ;
      RECT 61.55 53.23 61.83 53.51 ;
      RECT 61.55 53.03 61.71 53.51 ;
      RECT 60.73 53.03 61.71 53.19 ;
      RECT 60.73 50.98 60.89 53.19 ;
      RECT 60.69 52.54 60.89 52.82 ;
      RECT 60.35 50.98 60.89 51.14 ;
      RECT 60.35 50.8 60.57 51.14 ;
      RECT 60.25 56.67 60.41 61.86 ;
      RECT 60.25 56.67 61.69 56.83 ;
      RECT 61.53 56 61.69 56.83 ;
      RECT 60.41 54.4 60.57 56.83 ;
      RECT 61.39 26.36 61.55 26.72 ;
      RECT 59.25 26.36 61.55 26.52 ;
      RECT 59.25 26.04 59.41 26.52 ;
      RECT 58.6 26.04 59.41 26.2 ;
      RECT 61.37 50.66 61.53 51.5 ;
      RECT 60.73 50.66 61.53 50.82 ;
      RECT 60.73 50.18 60.89 50.82 ;
      RECT 60.25 50.18 60.89 50.5 ;
      RECT 60.25 47.07 60.41 50.5 ;
      RECT 60.25 47.07 60.73 47.23 ;
      RECT 60.57 45.44 60.73 47.23 ;
      RECT 61.13 55.68 61.29 56.51 ;
      RECT 61.13 55.68 61.53 55.84 ;
      RECT 61.37 53.67 61.53 55.84 ;
      RECT 60.89 53.67 61.53 53.83 ;
      RECT 60.89 53.35 61.17 53.83 ;
      RECT 61.37 62.9 61.53 67.89 ;
      RECT 61.31 65.82 61.53 66.55 ;
      RECT 61.05 51.7 61.43 51.92 ;
      RECT 61.05 50.98 61.21 51.92 ;
      RECT 59.22 28.01 61.38 28.17 ;
      RECT 61.22 27.34 61.38 28.17 ;
      RECT 61.06 27.93 61.38 28.17 ;
      RECT 60.22 26.97 60.38 28.17 ;
      RECT 59.22 26.68 59.38 28.17 ;
      RECT 60.57 47.39 60.73 49.72 ;
      RECT 60.57 47.39 61.05 47.55 ;
      RECT 60.89 43.85 61.05 47.55 ;
      RECT 60.27 43.85 61.05 44.01 ;
      RECT 60.27 39.56 60.43 44.01 ;
      RECT 60.27 39.56 60.61 39.84 ;
      RECT 60.45 39.16 60.61 39.84 ;
      RECT 60.73 24.79 60.93 25.35 ;
      RECT 60.61 24.79 60.93 25.03 ;
      RECT 60.59 34.44 60.93 34.72 ;
      RECT 60.77 32.44 60.93 34.72 ;
      RECT 60.59 33.11 60.93 33.39 ;
      RECT 60.59 32.44 60.93 32.72 ;
      RECT 60.59 40.7 60.93 40.98 ;
      RECT 60.77 38.7 60.93 40.98 ;
      RECT 60.59 40.03 60.93 40.31 ;
      RECT 60.59 38.7 60.93 38.98 ;
      RECT 60.61 21.85 60.77 24.3 ;
      RECT 60.61 21.85 60.91 22.13 ;
      RECT 60.73 54.06 60.89 56.51 ;
      RECT 60.37 54.06 60.89 54.22 ;
      RECT 60.37 52.98 60.57 54.22 ;
      RECT 60.37 51.34 60.53 54.22 ;
      RECT 60.37 51.34 60.57 52.12 ;
      RECT 60.43 12.56 60.59 13.61 ;
      RECT 60.53 11.9 60.69 13.24 ;
      RECT 59.41 11.9 60.69 12.06 ;
      RECT 60.35 9.6 60.51 12.06 ;
      RECT 59 18.3 59.94 18.46 ;
      RECT 59 17.05 59.36 18.46 ;
      RECT 59.2 16.2 59.36 18.46 ;
      RECT 59.15 16.2 60.11 16.36 ;
      RECT 59.88 16.07 60.55 16.23 ;
      RECT 59.15 16.08 59.31 16.36 ;
      RECT 60.19 8.96 60.51 9.12 ;
      RECT 60.35 7.8 60.51 9.12 ;
      RECT 58.01 7.91 58.17 8.8 ;
      RECT 58.01 7.91 59.09 8.07 ;
      RECT 58.93 7.8 60.51 7.96 ;
      RECT 59.52 16.52 59.7 16.84 ;
      RECT 59.52 16.52 60.42 16.68 ;
      RECT 59.93 46.75 60.09 47.43 ;
      RECT 59.61 46.75 60.41 46.91 ;
      RECT 60.25 44.23 60.41 46.91 ;
      RECT 59.61 44.23 59.77 46.91 ;
      RECT 60 16.92 60.16 18.12 ;
      RECT 60 16.92 60.4 17.08 ;
      RECT 58.85 11.5 59.01 13.22 ;
      RECT 58.85 12.22 60.37 12.38 ;
      RECT 58.85 11.5 59.27 11.66 ;
      RECT 59.77 26.02 60.33 26.18 ;
      RECT 59.77 25.58 59.93 26.18 ;
      RECT 59.23 25.58 59.93 25.74 ;
      RECT 59.23 24 59.43 25.74 ;
      RECT 58.43 24.3 59.43 24.46 ;
      RECT 59.23 22.71 59.39 25.74 ;
      RECT 59.33 22.04 59.49 22.99 ;
      RECT 59.49 21.85 59.65 22.32 ;
      RECT 58.81 22.13 59.17 22.41 ;
      RECT 59.01 21.53 59.17 22.41 ;
      RECT 59.88 21.53 60.04 21.92 ;
      RECT 59.01 21.53 60.04 21.69 ;
      RECT 59.7 20.21 59.86 21.69 ;
      RECT 59.74 26.69 59.9 27.85 ;
      RECT 59.7 26.69 59.94 27.33 ;
      RECT 57.71 34.88 59.91 35.04 ;
      RECT 59.63 34.59 59.91 35.04 ;
      RECT 58.69 34.59 58.93 35.04 ;
      RECT 57.71 34.59 57.99 35.04 ;
      RECT 58.69 38.38 58.93 39.02 ;
      RECT 59.63 38.38 59.91 38.83 ;
      RECT 57.71 38.38 57.99 38.83 ;
      RECT 57.71 38.38 59.91 38.54 ;
      RECT 59.55 23.18 59.71 23.84 ;
      RECT 59.55 23.18 59.88 23.34 ;
      RECT 59.72 22.65 59.88 23.34 ;
      RECT 57.87 36.47 59.75 36.63 ;
      RECT 59.59 35.86 59.75 36.63 ;
      RECT 58.73 35.23 58.89 36.63 ;
      RECT 57.87 35.86 58.03 36.63 ;
      RECT 59.69 35.23 59.85 36.05 ;
      RECT 57.77 35.23 57.93 36.05 ;
      RECT 59.69 37.11 59.85 38.19 ;
      RECT 58.73 36.79 58.89 38.19 ;
      RECT 57.77 37.11 57.93 38.19 ;
      RECT 59.59 36.79 59.75 37.39 ;
      RECT 57.87 36.79 58.03 37.39 ;
      RECT 57.87 36.79 59.75 36.95 ;
      RECT 58.49 50.66 58.65 51.5 ;
      RECT 58.49 50.66 59.29 50.82 ;
      RECT 59.13 50.18 59.29 50.82 ;
      RECT 59.13 50.18 59.77 50.5 ;
      RECT 59.61 47.07 59.77 50.5 ;
      RECT 59.29 47.07 59.77 47.23 ;
      RECT 59.29 45.44 59.45 47.23 ;
      RECT 59.61 56.67 59.77 61.86 ;
      RECT 58.33 56.67 59.77 56.83 ;
      RECT 59.45 54.4 59.61 56.83 ;
      RECT 58.33 56 58.49 56.83 ;
      RECT 59.29 47.39 59.45 49.72 ;
      RECT 58.97 47.39 59.45 47.55 ;
      RECT 58.97 43.85 59.13 47.55 ;
      RECT 58.97 43.85 59.75 44.01 ;
      RECT 59.59 39.56 59.75 44.01 ;
      RECT 59.41 39.56 59.75 39.84 ;
      RECT 59.41 39.16 59.57 39.84 ;
      RECT 58.2 28.52 59.29 28.68 ;
      RECT 59.01 28.35 59.29 28.68 ;
      RECT 59.01 28.35 59.69 28.51 ;
      RECT 58.19 53.23 58.47 53.51 ;
      RECT 58.31 53.03 58.47 53.51 ;
      RECT 58.31 53.03 59.29 53.19 ;
      RECT 59.13 50.98 59.29 53.19 ;
      RECT 59.13 52.54 59.33 52.82 ;
      RECT 59.13 50.98 59.67 51.14 ;
      RECT 59.45 50.8 59.67 51.14 ;
      RECT 57.85 68.07 59.67 68.23 ;
      RECT 59.51 62.02 59.67 68.23 ;
      RECT 59.29 62.02 59.67 62.18 ;
      RECT 59.29 57.45 59.45 62.18 ;
      RECT 57.85 57.45 59.45 57.61 ;
      RECT 57.85 57.39 58.17 57.61 ;
      RECT 58.01 53.74 58.17 57.61 ;
      RECT 57.85 51.32 58.01 53.9 ;
      RECT 57.85 51.32 58.33 51.48 ;
      RECT 58.17 49.88 58.33 51.48 ;
      RECT 58.17 49.88 58.65 50.04 ;
      RECT 58.49 47.71 58.65 50.04 ;
      RECT 58.49 47.71 59.11 47.99 ;
      RECT 59.13 54.06 59.29 56.51 ;
      RECT 59.13 54.06 59.65 54.22 ;
      RECT 59.49 51.34 59.65 54.22 ;
      RECT 59.45 52.98 59.65 54.22 ;
      RECT 59.45 51.34 59.65 52.12 ;
      RECT 58.33 12.92 58.49 13.67 ;
      RECT 58.33 12.92 58.69 13.08 ;
      RECT 58.53 9.68 58.69 13.08 ;
      RECT 58.49 9.68 58.69 11.89 ;
      RECT 58.49 9.68 59.47 9.84 ;
      RECT 59.31 8.6 59.47 9.84 ;
      RECT 59.09 34.44 59.43 34.72 ;
      RECT 59.09 32.44 59.25 34.72 ;
      RECT 59.09 33.11 59.43 33.39 ;
      RECT 59.09 32.44 59.43 32.72 ;
      RECT 59.09 40.7 59.43 40.98 ;
      RECT 59.09 38.7 59.25 40.98 ;
      RECT 59.09 40.03 59.43 40.31 ;
      RECT 59.09 38.7 59.43 38.98 ;
      RECT 58.73 55.68 58.89 56.51 ;
      RECT 58.49 55.68 58.89 55.84 ;
      RECT 58.49 53.67 58.65 55.84 ;
      RECT 58.49 53.67 59.13 53.83 ;
      RECT 58.85 53.35 59.13 53.83 ;
      RECT 58.68 16.52 58.84 18.9 ;
      RECT 58.68 16.52 59.04 16.8 ;
      RECT 58.81 15.31 58.97 16.8 ;
      RECT 58.28 24.79 58.44 28.32 ;
      RECT 58.28 25.16 58.97 25.32 ;
      RECT 58.59 51.7 58.97 51.92 ;
      RECT 58.81 50.98 58.97 51.92 ;
      RECT 58.17 52.58 58.93 52.86 ;
      RECT 58.77 52.18 58.93 52.86 ;
      RECT 58.17 51.64 58.33 52.86 ;
      RECT 58.01 23.98 58.19 24.52 ;
      RECT 58.01 23.98 58.71 24.14 ;
      RECT 58.55 23.27 58.71 24.14 ;
      RECT 58.49 21.78 58.65 23.43 ;
      RECT 58.63 21.21 58.79 21.94 ;
      RECT 58.76 20.95 58.92 21.37 ;
      RECT 57.53 7.5 57.69 8.72 ;
      RECT 57.53 7.58 57.74 7.9 ;
      RECT 57.53 7.59 58.77 7.75 ;
      RECT 57.53 7.58 57.81 7.75 ;
      RECT 58.49 62.9 58.65 67.89 ;
      RECT 58.49 65.82 58.71 66.55 ;
      RECT 58.17 47.39 58.33 49.72 ;
      RECT 58.17 47.39 58.65 47.55 ;
      RECT 58.49 43.85 58.65 47.55 ;
      RECT 57.87 43.85 58.65 44.01 ;
      RECT 57.87 39.56 58.03 44.01 ;
      RECT 57.87 39.56 58.21 39.84 ;
      RECT 58.05 39.16 58.21 39.84 ;
      RECT 58.19 34.44 58.53 34.72 ;
      RECT 58.37 32.44 58.53 34.72 ;
      RECT 58.19 33.11 58.53 33.39 ;
      RECT 58.19 32.44 58.53 32.72 ;
      RECT 58.19 40.7 58.53 40.98 ;
      RECT 58.37 38.7 58.53 40.98 ;
      RECT 58.19 40.03 58.53 40.31 ;
      RECT 58.19 38.7 58.53 38.98 ;
      RECT 57.76 15.57 57.92 17.28 ;
      RECT 58.36 16.43 58.52 16.71 ;
      RECT 57.76 16.43 58.52 16.59 ;
      RECT 57.7 15.57 57.98 15.73 ;
      RECT 58.2 17.18 58.36 18.9 ;
      RECT 57.53 17.96 58.36 18.12 ;
      RECT 57.53 17.84 57.69 18.12 ;
      RECT 58.24 17.06 58.4 17.34 ;
      RECT 57.85 23.66 58.39 23.82 ;
      RECT 57.85 20.12 58.01 23.82 ;
      RECT 57.85 23.22 58.31 23.38 ;
      RECT 57.76 20.83 58.01 21.11 ;
      RECT 57.85 20.12 58.28 20.28 ;
      RECT 58.01 62.9 58.17 67.89 ;
      RECT 58.01 64.59 58.29 65.31 ;
      RECT 58.05 10.08 58.21 11.89 ;
      RECT 57.47 10.08 58.21 10.24 ;
      RECT 57.53 8.88 57.69 10.24 ;
      RECT 57.53 46.75 57.69 47.43 ;
      RECT 57.21 46.75 58.01 46.91 ;
      RECT 57.85 44.23 58.01 46.91 ;
      RECT 57.21 44.23 57.37 46.91 ;
      RECT 57.8 26.15 57.96 28.96 ;
      RECT 57.77 26.15 57.96 26.51 ;
      RECT 55.31 34.88 57.51 35.04 ;
      RECT 57.23 34.59 57.51 35.04 ;
      RECT 56.29 34.59 56.53 35.04 ;
      RECT 55.31 34.59 55.59 35.04 ;
      RECT 56.29 38.38 56.53 39.02 ;
      RECT 57.23 38.38 57.51 38.83 ;
      RECT 55.31 38.38 55.59 38.83 ;
      RECT 55.31 38.38 57.51 38.54 ;
      RECT 55.47 36.47 57.35 36.63 ;
      RECT 57.19 35.88 57.35 36.63 ;
      RECT 56.33 35.23 56.49 36.63 ;
      RECT 55.47 35.88 55.63 36.63 ;
      RECT 57.29 35.23 57.45 36.06 ;
      RECT 55.37 35.23 55.53 36.06 ;
      RECT 57.29 37.11 57.45 38.19 ;
      RECT 56.33 36.79 56.49 38.19 ;
      RECT 55.37 37.11 55.53 38.19 ;
      RECT 57.19 36.79 57.35 37.39 ;
      RECT 55.47 36.79 55.63 37.39 ;
      RECT 55.47 36.79 57.35 36.95 ;
      RECT 55.55 68.07 57.37 68.23 ;
      RECT 55.55 62.02 55.71 68.23 ;
      RECT 55.55 62.02 55.93 62.18 ;
      RECT 55.77 57.45 55.93 62.18 ;
      RECT 55.77 57.45 57.37 57.61 ;
      RECT 57.05 57.39 57.37 57.61 ;
      RECT 57.05 53.74 57.21 57.61 ;
      RECT 57.21 51.32 57.37 53.9 ;
      RECT 56.89 51.32 57.37 51.48 ;
      RECT 56.89 49.88 57.05 51.48 ;
      RECT 56.57 49.88 57.05 50.04 ;
      RECT 56.57 47.71 56.73 50.04 ;
      RECT 56.11 47.71 56.73 47.99 ;
      RECT 56.89 47.39 57.05 49.72 ;
      RECT 56.57 47.39 57.05 47.55 ;
      RECT 56.57 43.85 56.73 47.55 ;
      RECT 56.57 43.85 57.35 44.01 ;
      RECT 57.19 39.56 57.35 44.01 ;
      RECT 57.01 39.56 57.35 39.84 ;
      RECT 57.01 39.16 57.17 39.84 ;
      RECT 57.05 62.9 57.21 67.89 ;
      RECT 56.93 64.59 57.21 65.31 ;
      RECT 56.29 52.58 57.05 52.86 ;
      RECT 56.89 51.64 57.05 52.86 ;
      RECT 56.29 52.18 56.45 52.86 ;
      RECT 56.69 34.44 57.03 34.72 ;
      RECT 56.69 32.44 56.85 34.72 ;
      RECT 56.69 33.11 57.03 33.39 ;
      RECT 56.69 32.44 57.03 32.72 ;
      RECT 56.69 40.7 57.03 40.98 ;
      RECT 56.69 38.7 56.85 40.98 ;
      RECT 56.69 40.03 57.03 40.31 ;
      RECT 56.69 38.7 57.03 38.98 ;
      RECT 56.75 53.23 57.03 53.51 ;
      RECT 56.75 53.03 56.91 53.51 ;
      RECT 55.93 53.03 56.91 53.19 ;
      RECT 55.93 50.98 56.09 53.19 ;
      RECT 55.89 52.54 56.09 52.82 ;
      RECT 55.55 50.98 56.09 51.14 ;
      RECT 55.55 50.8 55.77 51.14 ;
      RECT 55.45 56.67 55.61 61.86 ;
      RECT 55.45 56.67 56.89 56.83 ;
      RECT 56.73 56 56.89 56.83 ;
      RECT 55.61 54.4 55.77 56.83 ;
      RECT 48.89 12.95 56.73 13.55 ;
      RECT 56.13 8.34 56.73 13.55 ;
      RECT 48.89 8.34 49.49 13.55 ;
      RECT 48.89 8.34 56.73 8.88 ;
      RECT 48.89 26.87 56.73 27.47 ;
      RECT 56.13 18.71 56.73 27.47 ;
      RECT 48.89 18.71 49.49 27.47 ;
      RECT 48.89 24.41 56.73 25.01 ;
      RECT 48.89 18.71 56.73 19.31 ;
      RECT 56.57 50.66 56.73 51.5 ;
      RECT 55.93 50.66 56.73 50.82 ;
      RECT 55.93 50.18 56.09 50.82 ;
      RECT 55.45 50.18 56.09 50.5 ;
      RECT 55.45 47.07 55.61 50.5 ;
      RECT 55.45 47.07 55.93 47.23 ;
      RECT 55.77 45.44 55.93 47.23 ;
      RECT 56.33 55.68 56.49 56.51 ;
      RECT 56.33 55.68 56.73 55.84 ;
      RECT 56.57 53.67 56.73 55.84 ;
      RECT 56.09 53.67 56.73 53.83 ;
      RECT 56.09 53.35 56.37 53.83 ;
      RECT 56.57 62.9 56.73 67.89 ;
      RECT 56.51 65.82 56.73 66.55 ;
      RECT 56.25 51.7 56.63 51.92 ;
      RECT 56.25 50.98 56.41 51.92 ;
      RECT 55.77 47.39 55.93 49.72 ;
      RECT 55.77 47.39 56.25 47.55 ;
      RECT 56.09 43.85 56.25 47.55 ;
      RECT 55.47 43.85 56.25 44.01 ;
      RECT 55.47 39.56 55.63 44.01 ;
      RECT 55.47 39.56 55.81 39.84 ;
      RECT 55.65 39.16 55.81 39.84 ;
      RECT 55.79 34.44 56.13 34.72 ;
      RECT 55.97 32.44 56.13 34.72 ;
      RECT 55.79 33.11 56.13 33.39 ;
      RECT 55.79 32.44 56.13 32.72 ;
      RECT 55.79 40.7 56.13 40.98 ;
      RECT 55.97 38.7 56.13 40.98 ;
      RECT 55.79 40.03 56.13 40.31 ;
      RECT 55.79 38.7 56.13 38.98 ;
      RECT 55.93 54.06 56.09 56.51 ;
      RECT 55.57 54.06 56.09 54.22 ;
      RECT 55.57 52.98 55.77 54.22 ;
      RECT 55.57 51.34 55.73 54.22 ;
      RECT 55.57 51.34 55.77 52.12 ;
      RECT 55.13 46.75 55.29 47.43 ;
      RECT 54.81 46.75 55.61 46.91 ;
      RECT 55.45 44.23 55.61 46.91 ;
      RECT 54.81 44.23 54.97 46.91 ;
      RECT 52.91 34.88 55.11 35.04 ;
      RECT 54.83 34.59 55.11 35.04 ;
      RECT 53.89 34.59 54.13 35.04 ;
      RECT 52.91 34.59 53.19 35.04 ;
      RECT 53.89 38.38 54.13 39.02 ;
      RECT 54.83 38.38 55.11 38.83 ;
      RECT 52.91 38.38 53.19 38.83 ;
      RECT 52.91 38.38 55.11 38.54 ;
      RECT 53.07 36.47 54.95 36.63 ;
      RECT 54.79 35.86 54.95 36.63 ;
      RECT 53.93 35.23 54.09 36.63 ;
      RECT 53.07 35.86 53.23 36.63 ;
      RECT 54.89 35.23 55.05 36.05 ;
      RECT 52.97 35.23 53.13 36.05 ;
      RECT 54.89 37.11 55.05 38.19 ;
      RECT 53.93 36.79 54.09 38.19 ;
      RECT 52.97 37.11 53.13 38.19 ;
      RECT 54.79 36.79 54.95 37.39 ;
      RECT 53.07 36.79 53.23 37.39 ;
      RECT 53.07 36.79 54.95 36.95 ;
      RECT 53.69 50.66 53.85 51.5 ;
      RECT 53.69 50.66 54.49 50.82 ;
      RECT 54.33 50.18 54.49 50.82 ;
      RECT 54.33 50.18 54.97 50.5 ;
      RECT 54.81 47.07 54.97 50.5 ;
      RECT 54.49 47.07 54.97 47.23 ;
      RECT 54.49 45.44 54.65 47.23 ;
      RECT 54.81 56.67 54.97 61.86 ;
      RECT 53.53 56.67 54.97 56.83 ;
      RECT 54.65 54.4 54.81 56.83 ;
      RECT 53.53 56 53.69 56.83 ;
      RECT 54.49 47.39 54.65 49.72 ;
      RECT 54.17 47.39 54.65 47.55 ;
      RECT 54.17 43.85 54.33 47.55 ;
      RECT 54.17 43.85 54.95 44.01 ;
      RECT 54.79 39.56 54.95 44.01 ;
      RECT 54.61 39.56 54.95 39.84 ;
      RECT 54.61 39.16 54.77 39.84 ;
      RECT 53.39 53.23 53.67 53.51 ;
      RECT 53.51 53.03 53.67 53.51 ;
      RECT 53.51 53.03 54.49 53.19 ;
      RECT 54.33 50.98 54.49 53.19 ;
      RECT 54.33 52.54 54.53 52.82 ;
      RECT 54.33 50.98 54.87 51.14 ;
      RECT 54.65 50.8 54.87 51.14 ;
      RECT 53.05 68.07 54.87 68.23 ;
      RECT 54.71 62.02 54.87 68.23 ;
      RECT 54.49 62.02 54.87 62.18 ;
      RECT 54.49 57.45 54.65 62.18 ;
      RECT 53.05 57.45 54.65 57.61 ;
      RECT 53.05 57.39 53.37 57.61 ;
      RECT 53.21 53.74 53.37 57.61 ;
      RECT 53.05 51.32 53.21 53.9 ;
      RECT 53.05 51.32 53.53 51.48 ;
      RECT 53.37 49.88 53.53 51.48 ;
      RECT 53.37 49.88 53.85 50.04 ;
      RECT 53.69 47.71 53.85 50.04 ;
      RECT 53.69 47.71 54.31 47.99 ;
      RECT 54.33 54.06 54.49 56.51 ;
      RECT 54.33 54.06 54.85 54.22 ;
      RECT 54.69 51.34 54.85 54.22 ;
      RECT 54.65 52.98 54.85 54.22 ;
      RECT 54.65 51.34 54.85 52.12 ;
      RECT 54.29 34.44 54.63 34.72 ;
      RECT 54.29 32.44 54.45 34.72 ;
      RECT 54.29 33.11 54.63 33.39 ;
      RECT 54.29 32.44 54.63 32.72 ;
      RECT 54.29 40.7 54.63 40.98 ;
      RECT 54.29 38.7 54.45 40.98 ;
      RECT 54.29 40.03 54.63 40.31 ;
      RECT 54.29 38.7 54.63 38.98 ;
      RECT 53.93 55.68 54.09 56.51 ;
      RECT 53.69 55.68 54.09 55.84 ;
      RECT 53.69 53.67 53.85 55.84 ;
      RECT 53.69 53.67 54.33 53.83 ;
      RECT 54.05 53.35 54.33 53.83 ;
      RECT 53.79 51.7 54.17 51.92 ;
      RECT 54.01 50.98 54.17 51.92 ;
      RECT 53.37 52.58 54.13 52.86 ;
      RECT 53.97 52.18 54.13 52.86 ;
      RECT 53.37 51.64 53.53 52.86 ;
      RECT 53.69 62.9 53.85 67.89 ;
      RECT 53.69 65.82 53.91 66.55 ;
      RECT 53.37 47.39 53.53 49.72 ;
      RECT 53.37 47.39 53.85 47.55 ;
      RECT 53.69 43.85 53.85 47.55 ;
      RECT 53.07 43.85 53.85 44.01 ;
      RECT 53.07 39.56 53.23 44.01 ;
      RECT 53.07 39.56 53.41 39.84 ;
      RECT 53.25 39.16 53.41 39.84 ;
      RECT 53.39 34.44 53.73 34.72 ;
      RECT 53.57 32.44 53.73 34.72 ;
      RECT 53.39 33.11 53.73 33.39 ;
      RECT 53.39 32.44 53.73 32.72 ;
      RECT 53.39 40.7 53.73 40.98 ;
      RECT 53.57 38.7 53.73 40.98 ;
      RECT 53.39 40.03 53.73 40.31 ;
      RECT 53.39 38.7 53.73 38.98 ;
      RECT 53.21 62.9 53.37 67.89 ;
      RECT 53.21 64.59 53.49 65.31 ;
      RECT 52.73 46.75 52.89 47.43 ;
      RECT 52.41 46.75 53.21 46.91 ;
      RECT 53.05 44.23 53.21 46.91 ;
      RECT 52.41 44.23 52.57 46.91 ;
      RECT 50.51 34.88 52.71 35.04 ;
      RECT 52.43 34.59 52.71 35.04 ;
      RECT 51.49 34.59 51.73 35.04 ;
      RECT 50.51 34.59 50.79 35.04 ;
      RECT 51.49 38.38 51.73 39.02 ;
      RECT 52.43 38.38 52.71 38.83 ;
      RECT 50.51 38.38 50.79 38.83 ;
      RECT 50.51 38.38 52.71 38.54 ;
      RECT 50.67 36.47 52.55 36.63 ;
      RECT 52.39 35.88 52.55 36.63 ;
      RECT 51.53 35.23 51.69 36.63 ;
      RECT 50.67 35.88 50.83 36.63 ;
      RECT 52.49 35.23 52.65 36.06 ;
      RECT 50.57 35.23 50.73 36.06 ;
      RECT 52.49 37.11 52.65 38.19 ;
      RECT 51.53 36.79 51.69 38.19 ;
      RECT 50.57 37.11 50.73 38.19 ;
      RECT 52.39 36.79 52.55 37.39 ;
      RECT 50.67 36.79 50.83 37.39 ;
      RECT 50.67 36.79 52.55 36.95 ;
      RECT 50.75 68.07 52.57 68.23 ;
      RECT 50.75 62.02 50.91 68.23 ;
      RECT 50.75 62.02 51.13 62.18 ;
      RECT 50.97 57.45 51.13 62.18 ;
      RECT 50.97 57.45 52.57 57.61 ;
      RECT 52.25 57.39 52.57 57.61 ;
      RECT 52.25 53.74 52.41 57.61 ;
      RECT 52.41 51.32 52.57 53.9 ;
      RECT 52.09 51.32 52.57 51.48 ;
      RECT 52.09 49.88 52.25 51.48 ;
      RECT 51.77 49.88 52.25 50.04 ;
      RECT 51.77 47.71 51.93 50.04 ;
      RECT 51.31 47.71 51.93 47.99 ;
      RECT 52.09 47.39 52.25 49.72 ;
      RECT 51.77 47.39 52.25 47.55 ;
      RECT 51.77 43.85 51.93 47.55 ;
      RECT 51.77 43.85 52.55 44.01 ;
      RECT 52.39 39.56 52.55 44.01 ;
      RECT 52.21 39.56 52.55 39.84 ;
      RECT 52.21 39.16 52.37 39.84 ;
      RECT 52.25 62.9 52.41 67.89 ;
      RECT 52.13 64.59 52.41 65.31 ;
      RECT 51.49 52.58 52.25 52.86 ;
      RECT 52.09 51.64 52.25 52.86 ;
      RECT 51.49 52.18 51.65 52.86 ;
      RECT 51.89 34.44 52.23 34.72 ;
      RECT 51.89 32.44 52.05 34.72 ;
      RECT 51.89 33.11 52.23 33.39 ;
      RECT 51.89 32.44 52.23 32.72 ;
      RECT 51.89 40.7 52.23 40.98 ;
      RECT 51.89 38.7 52.05 40.98 ;
      RECT 51.89 40.03 52.23 40.31 ;
      RECT 51.89 38.7 52.23 38.98 ;
      RECT 51.95 53.23 52.23 53.51 ;
      RECT 51.95 53.03 52.11 53.51 ;
      RECT 51.13 53.03 52.11 53.19 ;
      RECT 51.13 50.98 51.29 53.19 ;
      RECT 51.09 52.54 51.29 52.82 ;
      RECT 50.75 50.98 51.29 51.14 ;
      RECT 50.75 50.8 50.97 51.14 ;
      RECT 50.65 56.67 50.81 61.86 ;
      RECT 50.65 56.67 52.09 56.83 ;
      RECT 51.93 56 52.09 56.83 ;
      RECT 50.81 54.4 50.97 56.83 ;
      RECT 51.77 50.66 51.93 51.5 ;
      RECT 51.13 50.66 51.93 50.82 ;
      RECT 51.13 50.18 51.29 50.82 ;
      RECT 50.65 50.18 51.29 50.5 ;
      RECT 50.65 47.07 50.81 50.5 ;
      RECT 50.65 47.07 51.13 47.23 ;
      RECT 50.97 45.44 51.13 47.23 ;
      RECT 51.53 55.68 51.69 56.51 ;
      RECT 51.53 55.68 51.93 55.84 ;
      RECT 51.77 53.67 51.93 55.84 ;
      RECT 51.29 53.67 51.93 53.83 ;
      RECT 51.29 53.35 51.57 53.83 ;
      RECT 51.77 62.9 51.93 67.89 ;
      RECT 51.71 65.82 51.93 66.55 ;
      RECT 51.45 51.7 51.83 51.92 ;
      RECT 51.45 50.98 51.61 51.92 ;
      RECT 50.97 47.39 51.13 49.72 ;
      RECT 50.97 47.39 51.45 47.55 ;
      RECT 51.29 43.85 51.45 47.55 ;
      RECT 50.67 43.85 51.45 44.01 ;
      RECT 50.67 39.56 50.83 44.01 ;
      RECT 50.67 39.56 51.01 39.84 ;
      RECT 50.85 39.16 51.01 39.84 ;
      RECT 50.99 34.44 51.33 34.72 ;
      RECT 51.17 32.44 51.33 34.72 ;
      RECT 50.99 33.11 51.33 33.39 ;
      RECT 50.99 32.44 51.33 32.72 ;
      RECT 50.99 40.7 51.33 40.98 ;
      RECT 51.17 38.7 51.33 40.98 ;
      RECT 50.99 40.03 51.33 40.31 ;
      RECT 50.99 38.7 51.33 38.98 ;
      RECT 51.13 54.06 51.29 56.51 ;
      RECT 50.77 54.06 51.29 54.22 ;
      RECT 50.77 52.98 50.97 54.22 ;
      RECT 50.77 51.34 50.93 54.22 ;
      RECT 50.77 51.34 50.97 52.12 ;
      RECT 50.33 46.75 50.49 47.43 ;
      RECT 50.01 46.75 50.81 46.91 ;
      RECT 50.65 44.23 50.81 46.91 ;
      RECT 50.01 44.23 50.17 46.91 ;
      RECT 48.11 34.88 50.31 35.04 ;
      RECT 50.03 34.59 50.31 35.04 ;
      RECT 49.09 34.59 49.33 35.04 ;
      RECT 48.11 34.59 48.39 35.04 ;
      RECT 49.09 38.38 49.33 39.02 ;
      RECT 50.03 38.38 50.31 38.83 ;
      RECT 48.11 38.38 48.39 38.83 ;
      RECT 48.11 38.38 50.31 38.54 ;
      RECT 48.27 36.47 50.15 36.63 ;
      RECT 49.99 35.86 50.15 36.63 ;
      RECT 49.13 35.23 49.29 36.63 ;
      RECT 48.27 35.86 48.43 36.63 ;
      RECT 50.09 35.23 50.25 36.05 ;
      RECT 48.17 35.23 48.33 36.05 ;
      RECT 50.09 37.11 50.25 38.19 ;
      RECT 49.13 36.79 49.29 38.19 ;
      RECT 48.17 37.11 48.33 38.19 ;
      RECT 49.99 36.79 50.15 37.39 ;
      RECT 48.27 36.79 48.43 37.39 ;
      RECT 48.27 36.79 50.15 36.95 ;
      RECT 48.89 50.66 49.05 51.5 ;
      RECT 48.89 50.66 49.69 50.82 ;
      RECT 49.53 50.18 49.69 50.82 ;
      RECT 49.53 50.18 50.17 50.5 ;
      RECT 50.01 47.07 50.17 50.5 ;
      RECT 49.69 47.07 50.17 47.23 ;
      RECT 49.69 45.44 49.85 47.23 ;
      RECT 50.01 56.67 50.17 61.86 ;
      RECT 48.73 56.67 50.17 56.83 ;
      RECT 49.85 54.4 50.01 56.83 ;
      RECT 48.73 56 48.89 56.83 ;
      RECT 49.69 47.39 49.85 49.72 ;
      RECT 49.37 47.39 49.85 47.55 ;
      RECT 49.37 43.85 49.53 47.55 ;
      RECT 49.37 43.85 50.15 44.01 ;
      RECT 49.99 39.56 50.15 44.01 ;
      RECT 49.81 39.56 50.15 39.84 ;
      RECT 49.81 39.16 49.97 39.84 ;
      RECT 48.59 53.23 48.87 53.51 ;
      RECT 48.71 53.03 48.87 53.51 ;
      RECT 48.71 53.03 49.69 53.19 ;
      RECT 49.53 50.98 49.69 53.19 ;
      RECT 49.53 52.54 49.73 52.82 ;
      RECT 49.53 50.98 50.07 51.14 ;
      RECT 49.85 50.8 50.07 51.14 ;
      RECT 48.25 68.07 50.07 68.23 ;
      RECT 49.91 62.02 50.07 68.23 ;
      RECT 49.69 62.02 50.07 62.18 ;
      RECT 49.69 57.45 49.85 62.18 ;
      RECT 48.25 57.45 49.85 57.61 ;
      RECT 48.25 57.39 48.57 57.61 ;
      RECT 48.41 53.74 48.57 57.61 ;
      RECT 48.25 51.32 48.41 53.9 ;
      RECT 48.25 51.32 48.73 51.48 ;
      RECT 48.57 49.88 48.73 51.48 ;
      RECT 48.57 49.88 49.05 50.04 ;
      RECT 48.89 47.71 49.05 50.04 ;
      RECT 48.89 47.71 49.51 47.99 ;
      RECT 49.53 54.06 49.69 56.51 ;
      RECT 49.53 54.06 50.05 54.22 ;
      RECT 49.89 51.34 50.05 54.22 ;
      RECT 49.85 52.98 50.05 54.22 ;
      RECT 49.85 51.34 50.05 52.12 ;
      RECT 49.49 34.44 49.83 34.72 ;
      RECT 49.49 32.44 49.65 34.72 ;
      RECT 49.49 33.11 49.83 33.39 ;
      RECT 49.49 32.44 49.83 32.72 ;
      RECT 49.49 40.7 49.83 40.98 ;
      RECT 49.49 38.7 49.65 40.98 ;
      RECT 49.49 40.03 49.83 40.31 ;
      RECT 49.49 38.7 49.83 38.98 ;
      RECT 49.13 55.68 49.29 56.51 ;
      RECT 48.89 55.68 49.29 55.84 ;
      RECT 48.89 53.67 49.05 55.84 ;
      RECT 48.89 53.67 49.53 53.83 ;
      RECT 49.25 53.35 49.53 53.83 ;
      RECT 48.99 51.7 49.37 51.92 ;
      RECT 49.21 50.98 49.37 51.92 ;
      RECT 48.57 52.58 49.33 52.86 ;
      RECT 49.17 52.18 49.33 52.86 ;
      RECT 48.57 51.64 48.73 52.86 ;
      RECT 48.89 62.9 49.05 67.89 ;
      RECT 48.89 65.82 49.11 66.55 ;
      RECT 48.57 47.39 48.73 49.72 ;
      RECT 48.57 47.39 49.05 47.55 ;
      RECT 48.89 43.85 49.05 47.55 ;
      RECT 48.27 43.85 49.05 44.01 ;
      RECT 48.27 39.56 48.43 44.01 ;
      RECT 48.27 39.56 48.61 39.84 ;
      RECT 48.45 39.16 48.61 39.84 ;
      RECT 46.61 6.84 48.21 7.24 ;
      RECT 47.61 6.24 49.01 6.84 ;
      RECT 45.81 6.24 47.21 6.84 ;
      RECT 48.59 34.44 48.93 34.72 ;
      RECT 48.77 32.44 48.93 34.72 ;
      RECT 48.59 33.11 48.93 33.39 ;
      RECT 48.59 32.44 48.93 32.72 ;
      RECT 48.59 40.7 48.93 40.98 ;
      RECT 48.77 38.7 48.93 40.98 ;
      RECT 48.59 40.03 48.93 40.31 ;
      RECT 48.59 38.7 48.93 38.98 ;
      RECT 48.41 62.9 48.57 67.89 ;
      RECT 48.41 64.59 48.69 65.31 ;
      RECT 47.93 46.75 48.09 47.43 ;
      RECT 47.93 46.75 48.41 46.91 ;
      RECT 48.25 44.23 48.41 46.91 ;
      RECT 46.73 46.75 46.89 47.43 ;
      RECT 46.41 46.75 46.89 46.91 ;
      RECT 46.41 44.23 46.57 46.91 ;
      RECT 44.51 34.88 46.71 35.04 ;
      RECT 46.43 34.59 46.71 35.04 ;
      RECT 45.49 34.59 45.73 35.04 ;
      RECT 44.51 34.59 44.79 35.04 ;
      RECT 45.49 38.38 45.73 39.02 ;
      RECT 46.43 38.38 46.71 38.83 ;
      RECT 44.51 38.38 44.79 38.83 ;
      RECT 44.51 38.38 46.71 38.54 ;
      RECT 44.67 36.47 46.55 36.63 ;
      RECT 46.39 35.88 46.55 36.63 ;
      RECT 45.53 35.23 45.69 36.63 ;
      RECT 44.67 35.88 44.83 36.63 ;
      RECT 46.49 35.23 46.65 36.06 ;
      RECT 44.57 35.23 44.73 36.06 ;
      RECT 46.49 37.11 46.65 38.19 ;
      RECT 45.53 36.79 45.69 38.19 ;
      RECT 44.57 37.11 44.73 38.19 ;
      RECT 46.39 36.79 46.55 37.39 ;
      RECT 44.67 36.79 44.83 37.39 ;
      RECT 44.67 36.79 46.55 36.95 ;
      RECT 44.75 68.07 46.57 68.23 ;
      RECT 44.75 62.02 44.91 68.23 ;
      RECT 44.75 62.02 45.13 62.18 ;
      RECT 44.97 57.45 45.13 62.18 ;
      RECT 44.97 57.45 46.57 57.61 ;
      RECT 46.25 57.39 46.57 57.61 ;
      RECT 46.25 53.74 46.41 57.61 ;
      RECT 46.41 51.32 46.57 53.9 ;
      RECT 46.09 51.32 46.57 51.48 ;
      RECT 46.09 49.88 46.25 51.48 ;
      RECT 45.77 49.88 46.25 50.04 ;
      RECT 45.77 47.71 45.93 50.04 ;
      RECT 45.31 47.71 45.93 47.99 ;
      RECT 46.09 47.39 46.25 49.72 ;
      RECT 45.77 47.39 46.25 47.55 ;
      RECT 45.77 43.85 45.93 47.55 ;
      RECT 45.77 43.85 46.55 44.01 ;
      RECT 46.39 39.56 46.55 44.01 ;
      RECT 46.21 39.56 46.55 39.84 ;
      RECT 46.21 39.16 46.37 39.84 ;
      RECT 46.25 62.9 46.41 67.89 ;
      RECT 46.13 64.59 46.41 65.31 ;
      RECT 45.49 52.58 46.25 52.86 ;
      RECT 46.09 51.64 46.25 52.86 ;
      RECT 45.49 52.18 45.65 52.86 ;
      RECT 45.89 34.44 46.23 34.72 ;
      RECT 45.89 32.44 46.05 34.72 ;
      RECT 45.89 33.11 46.23 33.39 ;
      RECT 45.89 32.44 46.23 32.72 ;
      RECT 45.89 40.7 46.23 40.98 ;
      RECT 45.89 38.7 46.05 40.98 ;
      RECT 45.89 40.03 46.23 40.31 ;
      RECT 45.89 38.7 46.23 38.98 ;
      RECT 45.95 53.23 46.23 53.51 ;
      RECT 45.95 53.03 46.11 53.51 ;
      RECT 45.13 53.03 46.11 53.19 ;
      RECT 45.13 50.98 45.29 53.19 ;
      RECT 45.09 52.54 45.29 52.82 ;
      RECT 44.75 50.98 45.29 51.14 ;
      RECT 44.75 50.8 44.97 51.14 ;
      RECT 44.65 56.67 44.81 61.86 ;
      RECT 44.65 56.67 46.09 56.83 ;
      RECT 45.93 56 46.09 56.83 ;
      RECT 44.81 54.4 44.97 56.83 ;
      RECT 38.09 12.95 45.93 13.55 ;
      RECT 45.33 8.34 45.93 13.55 ;
      RECT 38.09 8.34 38.69 13.55 ;
      RECT 38.09 8.34 45.93 8.88 ;
      RECT 38.09 26.87 45.93 27.47 ;
      RECT 45.33 18.71 45.93 27.47 ;
      RECT 38.09 18.71 38.69 27.47 ;
      RECT 38.09 24.41 45.93 25.01 ;
      RECT 38.09 18.71 45.93 19.31 ;
      RECT 45.77 50.66 45.93 51.5 ;
      RECT 45.13 50.66 45.93 50.82 ;
      RECT 45.13 50.18 45.29 50.82 ;
      RECT 44.65 50.18 45.29 50.5 ;
      RECT 44.65 47.07 44.81 50.5 ;
      RECT 44.65 47.07 45.13 47.23 ;
      RECT 44.97 45.44 45.13 47.23 ;
      RECT 45.53 55.68 45.69 56.51 ;
      RECT 45.53 55.68 45.93 55.84 ;
      RECT 45.77 53.67 45.93 55.84 ;
      RECT 45.29 53.67 45.93 53.83 ;
      RECT 45.29 53.35 45.57 53.83 ;
      RECT 45.77 62.9 45.93 67.89 ;
      RECT 45.71 65.82 45.93 66.55 ;
      RECT 45.45 51.7 45.83 51.92 ;
      RECT 45.45 50.98 45.61 51.92 ;
      RECT 44.97 47.39 45.13 49.72 ;
      RECT 44.97 47.39 45.45 47.55 ;
      RECT 45.29 43.85 45.45 47.55 ;
      RECT 44.67 43.85 45.45 44.01 ;
      RECT 44.67 39.56 44.83 44.01 ;
      RECT 44.67 39.56 45.01 39.84 ;
      RECT 44.85 39.16 45.01 39.84 ;
      RECT 44.99 34.44 45.33 34.72 ;
      RECT 45.17 32.44 45.33 34.72 ;
      RECT 44.99 33.11 45.33 33.39 ;
      RECT 44.99 32.44 45.33 32.72 ;
      RECT 44.99 40.7 45.33 40.98 ;
      RECT 45.17 38.7 45.33 40.98 ;
      RECT 44.99 40.03 45.33 40.31 ;
      RECT 44.99 38.7 45.33 38.98 ;
      RECT 45.13 54.06 45.29 56.51 ;
      RECT 44.77 54.06 45.29 54.22 ;
      RECT 44.77 52.98 44.97 54.22 ;
      RECT 44.77 51.34 44.93 54.22 ;
      RECT 44.77 51.34 44.97 52.12 ;
      RECT 44.33 46.75 44.49 47.43 ;
      RECT 44.01 46.75 44.81 46.91 ;
      RECT 44.65 44.23 44.81 46.91 ;
      RECT 44.01 44.23 44.17 46.91 ;
      RECT 42.11 34.88 44.31 35.04 ;
      RECT 44.03 34.59 44.31 35.04 ;
      RECT 43.09 34.59 43.33 35.04 ;
      RECT 42.11 34.59 42.39 35.04 ;
      RECT 43.09 38.38 43.33 39.02 ;
      RECT 44.03 38.38 44.31 38.83 ;
      RECT 42.11 38.38 42.39 38.83 ;
      RECT 42.11 38.38 44.31 38.54 ;
      RECT 42.27 36.47 44.15 36.63 ;
      RECT 43.99 35.86 44.15 36.63 ;
      RECT 43.13 35.23 43.29 36.63 ;
      RECT 42.27 35.86 42.43 36.63 ;
      RECT 44.09 35.23 44.25 36.05 ;
      RECT 42.17 35.23 42.33 36.05 ;
      RECT 44.09 37.11 44.25 38.19 ;
      RECT 43.13 36.79 43.29 38.19 ;
      RECT 42.17 37.11 42.33 38.19 ;
      RECT 43.99 36.79 44.15 37.39 ;
      RECT 42.27 36.79 42.43 37.39 ;
      RECT 42.27 36.79 44.15 36.95 ;
      RECT 42.89 50.66 43.05 51.5 ;
      RECT 42.89 50.66 43.69 50.82 ;
      RECT 43.53 50.18 43.69 50.82 ;
      RECT 43.53 50.18 44.17 50.5 ;
      RECT 44.01 47.07 44.17 50.5 ;
      RECT 43.69 47.07 44.17 47.23 ;
      RECT 43.69 45.44 43.85 47.23 ;
      RECT 44.01 56.67 44.17 61.86 ;
      RECT 42.73 56.67 44.17 56.83 ;
      RECT 43.85 54.4 44.01 56.83 ;
      RECT 42.73 56 42.89 56.83 ;
      RECT 43.69 47.39 43.85 49.72 ;
      RECT 43.37 47.39 43.85 47.55 ;
      RECT 43.37 43.85 43.53 47.55 ;
      RECT 43.37 43.85 44.15 44.01 ;
      RECT 43.99 39.56 44.15 44.01 ;
      RECT 43.81 39.56 44.15 39.84 ;
      RECT 43.81 39.16 43.97 39.84 ;
      RECT 42.59 53.23 42.87 53.51 ;
      RECT 42.71 53.03 42.87 53.51 ;
      RECT 42.71 53.03 43.69 53.19 ;
      RECT 43.53 50.98 43.69 53.19 ;
      RECT 43.53 52.54 43.73 52.82 ;
      RECT 43.53 50.98 44.07 51.14 ;
      RECT 43.85 50.8 44.07 51.14 ;
      RECT 42.25 68.07 44.07 68.23 ;
      RECT 43.91 62.02 44.07 68.23 ;
      RECT 43.69 62.02 44.07 62.18 ;
      RECT 43.69 57.45 43.85 62.18 ;
      RECT 42.25 57.45 43.85 57.61 ;
      RECT 42.25 57.39 42.57 57.61 ;
      RECT 42.41 53.74 42.57 57.61 ;
      RECT 42.25 51.32 42.41 53.9 ;
      RECT 42.25 51.32 42.73 51.48 ;
      RECT 42.57 49.88 42.73 51.48 ;
      RECT 42.57 49.88 43.05 50.04 ;
      RECT 42.89 47.71 43.05 50.04 ;
      RECT 42.89 47.71 43.51 47.99 ;
      RECT 43.53 54.06 43.69 56.51 ;
      RECT 43.53 54.06 44.05 54.22 ;
      RECT 43.89 51.34 44.05 54.22 ;
      RECT 43.85 52.98 44.05 54.22 ;
      RECT 43.85 51.34 44.05 52.12 ;
      RECT 43.49 34.44 43.83 34.72 ;
      RECT 43.49 32.44 43.65 34.72 ;
      RECT 43.49 33.11 43.83 33.39 ;
      RECT 43.49 32.44 43.83 32.72 ;
      RECT 43.49 40.7 43.83 40.98 ;
      RECT 43.49 38.7 43.65 40.98 ;
      RECT 43.49 40.03 43.83 40.31 ;
      RECT 43.49 38.7 43.83 38.98 ;
      RECT 43.13 55.68 43.29 56.51 ;
      RECT 42.89 55.68 43.29 55.84 ;
      RECT 42.89 53.67 43.05 55.84 ;
      RECT 42.89 53.67 43.53 53.83 ;
      RECT 43.25 53.35 43.53 53.83 ;
      RECT 42.99 51.7 43.37 51.92 ;
      RECT 43.21 50.98 43.37 51.92 ;
      RECT 42.57 52.58 43.33 52.86 ;
      RECT 43.17 52.18 43.33 52.86 ;
      RECT 42.57 51.64 42.73 52.86 ;
      RECT 42.89 62.9 43.05 67.89 ;
      RECT 42.89 65.82 43.11 66.55 ;
      RECT 42.57 47.39 42.73 49.72 ;
      RECT 42.57 47.39 43.05 47.55 ;
      RECT 42.89 43.85 43.05 47.55 ;
      RECT 42.27 43.85 43.05 44.01 ;
      RECT 42.27 39.56 42.43 44.01 ;
      RECT 42.27 39.56 42.61 39.84 ;
      RECT 42.45 39.16 42.61 39.84 ;
      RECT 42.59 34.44 42.93 34.72 ;
      RECT 42.77 32.44 42.93 34.72 ;
      RECT 42.59 33.11 42.93 33.39 ;
      RECT 42.59 32.44 42.93 32.72 ;
      RECT 42.59 40.7 42.93 40.98 ;
      RECT 42.77 38.7 42.93 40.98 ;
      RECT 42.59 40.03 42.93 40.31 ;
      RECT 42.59 38.7 42.93 38.98 ;
      RECT 42.41 62.9 42.57 67.89 ;
      RECT 42.41 64.59 42.69 65.31 ;
      RECT 41.93 46.75 42.09 47.43 ;
      RECT 41.61 46.75 42.41 46.91 ;
      RECT 42.25 44.23 42.41 46.91 ;
      RECT 41.61 44.23 41.77 46.91 ;
      RECT 39.71 34.88 41.91 35.04 ;
      RECT 41.63 34.59 41.91 35.04 ;
      RECT 40.69 34.59 40.93 35.04 ;
      RECT 39.71 34.59 39.99 35.04 ;
      RECT 40.69 38.38 40.93 39.02 ;
      RECT 41.63 38.38 41.91 38.83 ;
      RECT 39.71 38.38 39.99 38.83 ;
      RECT 39.71 38.38 41.91 38.54 ;
      RECT 39.87 36.47 41.75 36.63 ;
      RECT 41.59 35.88 41.75 36.63 ;
      RECT 40.73 35.23 40.89 36.63 ;
      RECT 39.87 35.88 40.03 36.63 ;
      RECT 41.69 35.23 41.85 36.06 ;
      RECT 39.77 35.23 39.93 36.06 ;
      RECT 41.69 37.11 41.85 38.19 ;
      RECT 40.73 36.79 40.89 38.19 ;
      RECT 39.77 37.11 39.93 38.19 ;
      RECT 41.59 36.79 41.75 37.39 ;
      RECT 39.87 36.79 40.03 37.39 ;
      RECT 39.87 36.79 41.75 36.95 ;
      RECT 39.95 68.07 41.77 68.23 ;
      RECT 39.95 62.02 40.11 68.23 ;
      RECT 39.95 62.02 40.33 62.18 ;
      RECT 40.17 57.45 40.33 62.18 ;
      RECT 40.17 57.45 41.77 57.61 ;
      RECT 41.45 57.39 41.77 57.61 ;
      RECT 41.45 53.74 41.61 57.61 ;
      RECT 41.61 51.32 41.77 53.9 ;
      RECT 41.29 51.32 41.77 51.48 ;
      RECT 41.29 49.88 41.45 51.48 ;
      RECT 40.97 49.88 41.45 50.04 ;
      RECT 40.97 47.71 41.13 50.04 ;
      RECT 40.51 47.71 41.13 47.99 ;
      RECT 41.29 47.39 41.45 49.72 ;
      RECT 40.97 47.39 41.45 47.55 ;
      RECT 40.97 43.85 41.13 47.55 ;
      RECT 40.97 43.85 41.75 44.01 ;
      RECT 41.59 39.56 41.75 44.01 ;
      RECT 41.41 39.56 41.75 39.84 ;
      RECT 41.41 39.16 41.57 39.84 ;
      RECT 41.45 62.9 41.61 67.89 ;
      RECT 41.33 64.59 41.61 65.31 ;
      RECT 40.69 52.58 41.45 52.86 ;
      RECT 41.29 51.64 41.45 52.86 ;
      RECT 40.69 52.18 40.85 52.86 ;
      RECT 41.09 34.44 41.43 34.72 ;
      RECT 41.09 32.44 41.25 34.72 ;
      RECT 41.09 33.11 41.43 33.39 ;
      RECT 41.09 32.44 41.43 32.72 ;
      RECT 41.09 40.7 41.43 40.98 ;
      RECT 41.09 38.7 41.25 40.98 ;
      RECT 41.09 40.03 41.43 40.31 ;
      RECT 41.09 38.7 41.43 38.98 ;
      RECT 41.15 53.23 41.43 53.51 ;
      RECT 41.15 53.03 41.31 53.51 ;
      RECT 40.33 53.03 41.31 53.19 ;
      RECT 40.33 50.98 40.49 53.19 ;
      RECT 40.29 52.54 40.49 52.82 ;
      RECT 39.95 50.98 40.49 51.14 ;
      RECT 39.95 50.8 40.17 51.14 ;
      RECT 39.85 56.67 40.01 61.86 ;
      RECT 39.85 56.67 41.29 56.83 ;
      RECT 41.13 56 41.29 56.83 ;
      RECT 40.01 54.4 40.17 56.83 ;
      RECT 40.97 50.66 41.13 51.5 ;
      RECT 40.33 50.66 41.13 50.82 ;
      RECT 40.33 50.18 40.49 50.82 ;
      RECT 39.85 50.18 40.49 50.5 ;
      RECT 39.85 47.07 40.01 50.5 ;
      RECT 39.85 47.07 40.33 47.23 ;
      RECT 40.17 45.44 40.33 47.23 ;
      RECT 40.73 55.68 40.89 56.51 ;
      RECT 40.73 55.68 41.13 55.84 ;
      RECT 40.97 53.67 41.13 55.84 ;
      RECT 40.49 53.67 41.13 53.83 ;
      RECT 40.49 53.35 40.77 53.83 ;
      RECT 40.97 62.9 41.13 67.89 ;
      RECT 40.91 65.82 41.13 66.55 ;
      RECT 40.65 51.7 41.03 51.92 ;
      RECT 40.65 50.98 40.81 51.92 ;
      RECT 40.17 47.39 40.33 49.72 ;
      RECT 40.17 47.39 40.65 47.55 ;
      RECT 40.49 43.85 40.65 47.55 ;
      RECT 39.87 43.85 40.65 44.01 ;
      RECT 39.87 39.56 40.03 44.01 ;
      RECT 39.87 39.56 40.21 39.84 ;
      RECT 40.05 39.16 40.21 39.84 ;
      RECT 40.19 34.44 40.53 34.72 ;
      RECT 40.37 32.44 40.53 34.72 ;
      RECT 40.19 33.11 40.53 33.39 ;
      RECT 40.19 32.44 40.53 32.72 ;
      RECT 40.19 40.7 40.53 40.98 ;
      RECT 40.37 38.7 40.53 40.98 ;
      RECT 40.19 40.03 40.53 40.31 ;
      RECT 40.19 38.7 40.53 38.98 ;
      RECT 40.33 54.06 40.49 56.51 ;
      RECT 39.97 54.06 40.49 54.22 ;
      RECT 39.97 52.98 40.17 54.22 ;
      RECT 39.97 51.34 40.13 54.22 ;
      RECT 39.97 51.34 40.17 52.12 ;
      RECT 39.53 46.75 39.69 47.43 ;
      RECT 39.21 46.75 40.01 46.91 ;
      RECT 39.85 44.23 40.01 46.91 ;
      RECT 39.21 44.23 39.37 46.91 ;
      RECT 37.31 34.88 39.51 35.04 ;
      RECT 39.23 34.59 39.51 35.04 ;
      RECT 38.29 34.59 38.53 35.04 ;
      RECT 37.31 34.59 37.59 35.04 ;
      RECT 38.29 38.38 38.53 39.02 ;
      RECT 39.23 38.38 39.51 38.83 ;
      RECT 37.31 38.38 37.59 38.83 ;
      RECT 37.31 38.38 39.51 38.54 ;
      RECT 37.47 36.47 39.35 36.63 ;
      RECT 39.19 35.86 39.35 36.63 ;
      RECT 38.33 35.23 38.49 36.63 ;
      RECT 37.47 35.86 37.63 36.63 ;
      RECT 39.29 35.23 39.45 36.05 ;
      RECT 37.37 35.23 37.53 36.05 ;
      RECT 39.29 37.11 39.45 38.19 ;
      RECT 38.33 36.79 38.49 38.19 ;
      RECT 37.37 37.11 37.53 38.19 ;
      RECT 39.19 36.79 39.35 37.39 ;
      RECT 37.47 36.79 37.63 37.39 ;
      RECT 37.47 36.79 39.35 36.95 ;
      RECT 38.09 50.66 38.25 51.5 ;
      RECT 38.09 50.66 38.89 50.82 ;
      RECT 38.73 50.18 38.89 50.82 ;
      RECT 38.73 50.18 39.37 50.5 ;
      RECT 39.21 47.07 39.37 50.5 ;
      RECT 38.89 47.07 39.37 47.23 ;
      RECT 38.89 45.44 39.05 47.23 ;
      RECT 39.21 56.67 39.37 61.86 ;
      RECT 37.93 56.67 39.37 56.83 ;
      RECT 39.05 54.4 39.21 56.83 ;
      RECT 37.93 56 38.09 56.83 ;
      RECT 38.89 47.39 39.05 49.72 ;
      RECT 38.57 47.39 39.05 47.55 ;
      RECT 38.57 43.85 38.73 47.55 ;
      RECT 38.57 43.85 39.35 44.01 ;
      RECT 39.19 39.56 39.35 44.01 ;
      RECT 39.01 39.56 39.35 39.84 ;
      RECT 39.01 39.16 39.17 39.84 ;
      RECT 37.79 53.23 38.07 53.51 ;
      RECT 37.91 53.03 38.07 53.51 ;
      RECT 37.91 53.03 38.89 53.19 ;
      RECT 38.73 50.98 38.89 53.19 ;
      RECT 38.73 52.54 38.93 52.82 ;
      RECT 38.73 50.98 39.27 51.14 ;
      RECT 39.05 50.8 39.27 51.14 ;
      RECT 37.45 68.07 39.27 68.23 ;
      RECT 39.11 62.02 39.27 68.23 ;
      RECT 38.89 62.02 39.27 62.18 ;
      RECT 38.89 57.45 39.05 62.18 ;
      RECT 37.45 57.45 39.05 57.61 ;
      RECT 37.45 57.39 37.77 57.61 ;
      RECT 37.61 53.74 37.77 57.61 ;
      RECT 37.45 51.32 37.61 53.9 ;
      RECT 37.45 51.32 37.93 51.48 ;
      RECT 37.77 49.88 37.93 51.48 ;
      RECT 37.77 49.88 38.25 50.04 ;
      RECT 38.09 47.71 38.25 50.04 ;
      RECT 38.09 47.71 38.71 47.99 ;
      RECT 38.73 54.06 38.89 56.51 ;
      RECT 38.73 54.06 39.25 54.22 ;
      RECT 39.09 51.34 39.25 54.22 ;
      RECT 39.05 52.98 39.25 54.22 ;
      RECT 39.05 51.34 39.25 52.12 ;
      RECT 38.69 34.44 39.03 34.72 ;
      RECT 38.69 32.44 38.85 34.72 ;
      RECT 38.69 33.11 39.03 33.39 ;
      RECT 38.69 32.44 39.03 32.72 ;
      RECT 38.69 40.7 39.03 40.98 ;
      RECT 38.69 38.7 38.85 40.98 ;
      RECT 38.69 40.03 39.03 40.31 ;
      RECT 38.69 38.7 39.03 38.98 ;
      RECT 38.33 55.68 38.49 56.51 ;
      RECT 38.09 55.68 38.49 55.84 ;
      RECT 38.09 53.67 38.25 55.84 ;
      RECT 38.09 53.67 38.73 53.83 ;
      RECT 38.45 53.35 38.73 53.83 ;
      RECT 38.19 51.7 38.57 51.92 ;
      RECT 38.41 50.98 38.57 51.92 ;
      RECT 37.77 52.58 38.53 52.86 ;
      RECT 38.37 52.18 38.53 52.86 ;
      RECT 37.77 51.64 37.93 52.86 ;
      RECT 38.09 62.9 38.25 67.89 ;
      RECT 38.09 65.82 38.31 66.55 ;
      RECT 37.77 47.39 37.93 49.72 ;
      RECT 37.77 47.39 38.25 47.55 ;
      RECT 38.09 43.85 38.25 47.55 ;
      RECT 37.47 43.85 38.25 44.01 ;
      RECT 37.47 39.56 37.63 44.01 ;
      RECT 37.47 39.56 37.81 39.84 ;
      RECT 37.65 39.16 37.81 39.84 ;
      RECT 37.79 34.44 38.13 34.72 ;
      RECT 37.97 32.44 38.13 34.72 ;
      RECT 37.79 33.11 38.13 33.39 ;
      RECT 37.79 32.44 38.13 32.72 ;
      RECT 37.79 40.7 38.13 40.98 ;
      RECT 37.97 38.7 38.13 40.98 ;
      RECT 37.79 40.03 38.13 40.31 ;
      RECT 37.79 38.7 38.13 38.98 ;
      RECT 37.61 62.9 37.77 67.89 ;
      RECT 37.61 64.59 37.89 65.31 ;
      RECT 37.13 46.75 37.29 47.43 ;
      RECT 36.81 46.75 37.61 46.91 ;
      RECT 37.45 44.23 37.61 46.91 ;
      RECT 36.81 44.23 36.97 46.91 ;
      RECT 36.61 10.08 36.77 11.89 ;
      RECT 36.61 10.08 37.35 10.24 ;
      RECT 37.13 8.88 37.29 10.24 ;
      RECT 37.13 7.5 37.29 8.72 ;
      RECT 37.08 7.58 37.29 7.9 ;
      RECT 36.05 7.59 37.29 7.75 ;
      RECT 37.01 7.58 37.29 7.75 ;
      RECT 29.09 15.8 29.25 16.08 ;
      RECT 25.97 15.8 26.13 16.08 ;
      RECT 28.49 15.8 29.25 15.96 ;
      RECT 25.97 15.8 26.73 15.96 ;
      RECT 26.57 14.07 26.73 15.96 ;
      RECT 34.99 14.25 35.15 15.89 ;
      RECT 20.07 14.25 20.23 15.89 ;
      RECT 27.53 12.21 27.69 15.8 ;
      RECT 28.49 14.07 28.65 15.96 ;
      RECT 32.47 14.12 32.65 15.79 ;
      RECT 31.19 14.1 31.35 15.79 ;
      RECT 23.87 14.1 24.03 15.79 ;
      RECT 22.57 14.12 22.75 15.79 ;
      RECT 36.33 14.64 36.49 15.6 ;
      RECT 18.73 14.64 18.89 15.6 ;
      RECT 37.13 12.64 37.29 14.96 ;
      RECT 17.93 12.64 18.09 14.96 ;
      RECT 30.15 14.1 30.31 14.89 ;
      RECT 24.91 14.1 25.07 14.89 ;
      RECT 34.71 14.64 37.29 14.84 ;
      RECT 17.93 14.64 20.51 14.84 ;
      RECT 20.35 12.56 20.51 14.84 ;
      RECT 34.71 14.25 36.16 14.84 ;
      RECT 19.06 14.25 20.51 14.84 ;
      RECT 29.21 14.36 30.31 14.52 ;
      RECT 24.91 14.36 26.01 14.52 ;
      RECT 25.85 14.08 26.01 14.52 ;
      RECT 29.21 14.08 29.37 14.52 ;
      RECT 31.19 14.12 34.87 14.28 ;
      RECT 19.06 14.25 24.03 14.28 ;
      RECT 30.15 14.1 31.67 14.26 ;
      RECT 23.55 14.1 25.07 14.26 ;
      RECT 20.35 14.12 25.07 14.26 ;
      RECT 28.49 14.08 29.37 14.24 ;
      RECT 25.85 14.08 26.73 14.24 ;
      RECT 26.39 14.07 28.83 14.23 ;
      RECT 34.71 12.56 34.87 14.84 ;
      RECT 33.75 12.55 33.91 14.28 ;
      RECT 32.87 13.45 33.03 14.28 ;
      RECT 22.19 13.45 22.35 14.28 ;
      RECT 21.31 12.55 21.47 14.28 ;
      RECT 30.41 12.32 30.57 14.26 ;
      RECT 24.65 12.32 24.81 14.26 ;
      RECT 28.67 13.38 28.83 14.24 ;
      RECT 26.39 13.38 26.55 14.24 ;
      RECT 32.79 12.55 32.95 13.61 ;
      RECT 22.27 12.55 22.43 13.61 ;
      RECT 28.55 13.38 28.83 13.54 ;
      RECT 26.39 13.38 26.67 13.54 ;
      RECT 36.46 17.18 36.62 18.9 ;
      RECT 36.46 17.96 37.29 18.12 ;
      RECT 37.13 17.84 37.29 18.12 ;
      RECT 36.42 17.06 36.58 17.34 ;
      RECT 35.44 19.61 35.6 21.25 ;
      RECT 28.49 20.42 28.65 21.25 ;
      RECT 27.53 16.39 27.69 21.25 ;
      RECT 26.57 20.42 26.73 21.25 ;
      RECT 19.62 19.61 19.78 21.25 ;
      RECT 36.22 20.89 36.64 21.05 ;
      RECT 34.48 19.61 34.64 21.05 ;
      RECT 20.58 19.61 20.74 21.05 ;
      RECT 18.58 20.89 19 21.05 ;
      RECT 18.84 19.61 19 21.05 ;
      RECT 33.48 20.21 33.64 20.89 ;
      RECT 31.23 20.43 31.39 20.89 ;
      RECT 23.83 20.43 23.99 20.89 ;
      RECT 21.58 20.21 21.74 20.89 ;
      RECT 36.22 19.61 36.38 21.05 ;
      RECT 30.77 20.43 31.39 20.59 ;
      RECT 23.83 20.43 24.45 20.59 ;
      RECT 24.29 19.1 24.45 20.59 ;
      RECT 28.57 19.16 28.73 20.58 ;
      RECT 26.49 19.16 26.65 20.58 ;
      RECT 29.81 19.16 29.97 20.49 ;
      RECT 25.25 19.16 25.41 20.49 ;
      RECT 30.77 19.1 30.93 20.59 ;
      RECT 33.48 20.21 34.64 20.37 ;
      RECT 34.44 19.61 34.64 20.37 ;
      RECT 20.58 20.21 21.74 20.37 ;
      RECT 20.58 19.61 20.78 20.37 ;
      RECT 34.44 19.61 35.6 19.81 ;
      RECT 19.62 19.61 20.78 19.81 ;
      RECT 34.27 19.61 37.21 19.77 ;
      RECT 18.01 19.61 20.95 19.77 ;
      RECT 20.79 19.1 20.95 19.77 ;
      RECT 33.31 19.1 33.59 19.73 ;
      RECT 21.63 19.1 21.91 19.73 ;
      RECT 34.27 19.1 34.43 19.77 ;
      RECT 29.81 19.16 30.93 19.37 ;
      RECT 24.29 19.16 25.41 19.37 ;
      RECT 24.29 19.16 30.93 19.32 ;
      RECT 29.92 19.1 34.43 19.26 ;
      RECT 29.45 18.46 29.61 19.32 ;
      RECT 28.49 17.56 28.65 19.32 ;
      RECT 26.57 17.56 26.73 19.32 ;
      RECT 25.61 18.46 25.77 19.32 ;
      RECT 20.79 19.1 25.3 19.26 ;
      RECT 24.16 17.76 24.32 19.26 ;
      RECT 30.9 19.01 32.82 19.26 ;
      RECT 32.64 16.65 32.82 19.26 ;
      RECT 22.4 19.01 24.32 19.26 ;
      RECT 31.7 17.58 31.86 19.26 ;
      RECT 30.9 17.76 31.06 19.26 ;
      RECT 23.36 17.58 23.52 19.26 ;
      RECT 22.4 16.65 22.58 19.26 ;
      RECT 30.37 17.76 31.06 17.92 ;
      RECT 24.16 17.76 24.85 17.92 ;
      RECT 24.69 16.77 24.85 17.92 ;
      RECT 30.37 16.77 30.53 17.92 ;
      RECT 36.9 15.57 37.06 17.28 ;
      RECT 36.3 16.43 36.46 16.71 ;
      RECT 36.3 16.43 37.06 16.59 ;
      RECT 36.84 15.57 37.12 15.73 ;
      RECT 34.91 34.88 37.11 35.04 ;
      RECT 36.83 34.59 37.11 35.04 ;
      RECT 35.89 34.59 36.13 35.04 ;
      RECT 34.91 34.59 35.19 35.04 ;
      RECT 35.89 38.38 36.13 39.02 ;
      RECT 36.83 38.38 37.11 38.83 ;
      RECT 34.91 38.38 35.19 38.83 ;
      RECT 34.91 38.38 37.11 38.54 ;
      RECT 36.43 23.66 36.97 23.82 ;
      RECT 36.81 20.12 36.97 23.82 ;
      RECT 36.51 23.22 36.97 23.38 ;
      RECT 36.81 20.83 37.06 21.11 ;
      RECT 36.54 20.12 36.97 20.28 ;
      RECT 36.86 26.15 37.02 28.96 ;
      RECT 36.86 26.15 37.05 26.51 ;
      RECT 35.07 36.47 36.95 36.63 ;
      RECT 36.79 35.88 36.95 36.63 ;
      RECT 35.93 35.23 36.09 36.63 ;
      RECT 35.07 35.88 35.23 36.63 ;
      RECT 36.89 35.23 37.05 36.06 ;
      RECT 34.97 35.23 35.13 36.06 ;
      RECT 36.89 37.11 37.05 38.19 ;
      RECT 35.93 36.79 36.09 38.19 ;
      RECT 34.97 37.11 35.13 38.19 ;
      RECT 36.79 36.79 36.95 37.39 ;
      RECT 35.07 36.79 35.23 37.39 ;
      RECT 35.07 36.79 36.95 36.95 ;
      RECT 35.15 68.07 36.97 68.23 ;
      RECT 35.15 62.02 35.31 68.23 ;
      RECT 35.15 62.02 35.53 62.18 ;
      RECT 35.37 57.45 35.53 62.18 ;
      RECT 35.37 57.45 36.97 57.61 ;
      RECT 36.65 57.39 36.97 57.61 ;
      RECT 36.65 53.74 36.81 57.61 ;
      RECT 36.81 51.32 36.97 53.9 ;
      RECT 36.49 51.32 36.97 51.48 ;
      RECT 36.49 49.88 36.65 51.48 ;
      RECT 36.17 49.88 36.65 50.04 ;
      RECT 36.17 47.71 36.33 50.04 ;
      RECT 35.71 47.71 36.33 47.99 ;
      RECT 36.49 47.39 36.65 49.72 ;
      RECT 36.17 47.39 36.65 47.55 ;
      RECT 36.17 43.85 36.33 47.55 ;
      RECT 36.17 43.85 36.95 44.01 ;
      RECT 36.79 39.56 36.95 44.01 ;
      RECT 36.61 39.56 36.95 39.84 ;
      RECT 36.61 39.16 36.77 39.84 ;
      RECT 34.31 8.96 34.63 9.12 ;
      RECT 34.31 7.8 34.47 9.12 ;
      RECT 36.65 7.91 36.81 8.8 ;
      RECT 35.73 7.91 36.81 8.07 ;
      RECT 34.31 7.8 35.89 7.96 ;
      RECT 36.63 23.98 36.81 24.52 ;
      RECT 36.11 23.98 36.81 24.14 ;
      RECT 36.11 23.27 36.27 24.14 ;
      RECT 36.17 21.78 36.33 23.43 ;
      RECT 36.03 21.21 36.19 21.94 ;
      RECT 35.9 20.95 36.06 21.37 ;
      RECT 36.65 62.9 36.81 67.89 ;
      RECT 36.53 64.59 36.81 65.31 ;
      RECT 35.89 52.58 36.65 52.86 ;
      RECT 36.49 51.64 36.65 52.86 ;
      RECT 35.89 52.18 36.05 52.86 ;
      RECT 36.29 34.44 36.63 34.72 ;
      RECT 36.29 32.44 36.45 34.72 ;
      RECT 36.29 33.11 36.63 33.39 ;
      RECT 36.29 32.44 36.63 32.72 ;
      RECT 36.29 40.7 36.63 40.98 ;
      RECT 36.29 38.7 36.45 40.98 ;
      RECT 36.29 40.03 36.63 40.31 ;
      RECT 36.29 38.7 36.63 38.98 ;
      RECT 36.35 53.23 36.63 53.51 ;
      RECT 36.35 53.03 36.51 53.51 ;
      RECT 35.53 53.03 36.51 53.19 ;
      RECT 35.53 50.98 35.69 53.19 ;
      RECT 35.49 52.54 35.69 52.82 ;
      RECT 35.15 50.98 35.69 51.14 ;
      RECT 35.15 50.8 35.37 51.14 ;
      RECT 35.53 28.52 36.62 28.68 ;
      RECT 35.53 28.35 35.81 28.68 ;
      RECT 35.13 28.35 35.81 28.51 ;
      RECT 36.38 24.79 36.54 28.32 ;
      RECT 35.85 25.16 36.54 25.32 ;
      RECT 36.33 12.92 36.49 13.67 ;
      RECT 36.13 12.92 36.49 13.08 ;
      RECT 36.13 9.68 36.29 13.08 ;
      RECT 36.13 9.68 36.33 11.89 ;
      RECT 35.35 9.68 36.33 9.84 ;
      RECT 35.35 8.6 35.51 9.84 ;
      RECT 35.05 56.67 35.21 61.86 ;
      RECT 35.05 56.67 36.49 56.83 ;
      RECT 36.33 56 36.49 56.83 ;
      RECT 35.21 54.4 35.37 56.83 ;
      RECT 34.49 26.02 35.05 26.18 ;
      RECT 34.89 25.58 35.05 26.18 ;
      RECT 34.89 25.58 35.59 25.74 ;
      RECT 35.43 22.71 35.59 25.74 ;
      RECT 35.39 24 35.59 25.74 ;
      RECT 35.39 24.3 36.39 24.46 ;
      RECT 35.33 22.04 35.49 22.99 ;
      RECT 35.17 21.85 35.33 22.32 ;
      RECT 36.17 50.66 36.33 51.5 ;
      RECT 35.53 50.66 36.33 50.82 ;
      RECT 35.53 50.18 35.69 50.82 ;
      RECT 35.05 50.18 35.69 50.5 ;
      RECT 35.05 47.07 35.21 50.5 ;
      RECT 35.05 47.07 35.53 47.23 ;
      RECT 35.37 45.44 35.53 47.23 ;
      RECT 35.93 55.68 36.09 56.51 ;
      RECT 35.93 55.68 36.33 55.84 ;
      RECT 36.17 53.67 36.33 55.84 ;
      RECT 35.69 53.67 36.33 53.83 ;
      RECT 35.69 53.35 35.97 53.83 ;
      RECT 36.17 62.9 36.33 67.89 ;
      RECT 36.11 65.82 36.33 66.55 ;
      RECT 35.85 51.7 36.23 51.92 ;
      RECT 35.85 50.98 36.01 51.92 ;
      RECT 33.27 26.36 33.43 26.72 ;
      RECT 33.27 26.36 35.57 26.52 ;
      RECT 35.41 26.04 35.57 26.52 ;
      RECT 35.41 26.04 36.22 26.2 ;
      RECT 35.98 16.52 36.14 18.9 ;
      RECT 35.78 16.52 36.14 16.8 ;
      RECT 35.85 15.31 36.01 16.8 ;
      RECT 35.65 22.13 36.01 22.41 ;
      RECT 35.65 21.53 35.81 22.41 ;
      RECT 34.78 21.53 34.94 21.92 ;
      RECT 34.78 21.53 35.81 21.69 ;
      RECT 34.96 20.21 35.12 21.69 ;
      RECT 35.81 11.5 35.97 13.22 ;
      RECT 34.45 12.22 35.97 12.38 ;
      RECT 35.55 11.5 35.97 11.66 ;
      RECT 35.37 47.39 35.53 49.72 ;
      RECT 35.37 47.39 35.85 47.55 ;
      RECT 35.69 43.85 35.85 47.55 ;
      RECT 35.07 43.85 35.85 44.01 ;
      RECT 35.07 39.56 35.23 44.01 ;
      RECT 35.07 39.56 35.41 39.84 ;
      RECT 35.25 39.16 35.41 39.84 ;
      RECT 34.88 18.3 35.82 18.46 ;
      RECT 35.46 17.05 35.82 18.46 ;
      RECT 35.46 16.2 35.62 18.46 ;
      RECT 34.71 16.2 35.67 16.36 ;
      RECT 35.51 16.08 35.67 16.36 ;
      RECT 34.27 16.07 34.94 16.23 ;
      RECT 35.39 34.44 35.73 34.72 ;
      RECT 35.57 32.44 35.73 34.72 ;
      RECT 35.39 33.11 35.73 33.39 ;
      RECT 35.39 32.44 35.73 32.72 ;
      RECT 35.39 40.7 35.73 40.98 ;
      RECT 35.57 38.7 35.73 40.98 ;
      RECT 35.39 40.03 35.73 40.31 ;
      RECT 35.39 38.7 35.73 38.98 ;
      RECT 35.53 54.06 35.69 56.51 ;
      RECT 35.17 54.06 35.69 54.22 ;
      RECT 35.17 52.98 35.37 54.22 ;
      RECT 35.17 51.34 35.33 54.22 ;
      RECT 35.17 51.34 35.37 52.12 ;
      RECT 33.44 28.01 35.6 28.17 ;
      RECT 35.44 26.68 35.6 28.17 ;
      RECT 34.44 26.97 34.6 28.17 ;
      RECT 33.44 27.93 33.76 28.17 ;
      RECT 33.44 27.34 33.6 28.17 ;
      RECT 34.23 12.56 34.39 13.61 ;
      RECT 34.13 11.9 34.29 13.24 ;
      RECT 34.13 11.9 35.41 12.06 ;
      RECT 34.31 9.6 34.47 12.06 ;
      RECT 35.12 16.52 35.3 16.84 ;
      RECT 34.4 16.52 35.3 16.68 ;
      RECT 35.11 23.18 35.27 23.84 ;
      RECT 34.94 23.18 35.27 23.34 ;
      RECT 34.94 22.65 35.1 23.34 ;
      RECT 34.73 46.75 34.89 47.43 ;
      RECT 34.41 46.75 35.21 46.91 ;
      RECT 35.05 44.23 35.21 46.91 ;
      RECT 34.41 44.23 34.57 46.91 ;
      RECT 34.92 26.69 35.08 27.85 ;
      RECT 34.88 26.69 35.12 27.33 ;
      RECT 34.79 9.28 34.95 11.72 ;
      RECT 33.83 8.12 33.99 11.72 ;
      RECT 32.87 8.5 33.03 11.72 ;
      RECT 31.21 9.63 31.37 11.4 ;
      RECT 31.21 9.95 33.03 10.11 ;
      RECT 31.9 9.79 32.06 10.11 ;
      RECT 34.83 8.12 35.03 9.84 ;
      RECT 31.15 9.63 31.66 9.79 ;
      RECT 33.83 9.28 35.03 9.44 ;
      RECT 32.83 8.5 33.14 8.78 ;
      RECT 32.83 8.56 33.99 8.72 ;
      RECT 29.85 28.74 34.97 28.9 ;
      RECT 33.05 27.92 33.21 28.9 ;
      RECT 31.61 27.92 31.77 28.9 ;
      RECT 34.66 16.92 34.82 18.12 ;
      RECT 34.42 16.92 34.82 17.08 ;
      RECT 32.51 34.88 34.71 35.04 ;
      RECT 34.43 34.59 34.71 35.04 ;
      RECT 33.49 34.59 33.73 35.04 ;
      RECT 32.51 34.59 32.79 35.04 ;
      RECT 33.49 38.38 33.73 39.02 ;
      RECT 34.43 38.38 34.71 38.83 ;
      RECT 32.51 38.38 32.79 38.83 ;
      RECT 32.51 38.38 34.71 38.54 ;
      RECT 32.33 21.69 32.49 26.21 ;
      RECT 33.57 24.34 33.73 26.2 ;
      RECT 31.09 24.35 31.25 26.2 ;
      RECT 34.45 24.04 34.67 25.52 ;
      RECT 30.15 24.04 30.37 25.52 ;
      RECT 33.57 24.46 34.67 24.63 ;
      RECT 30.15 24.46 31.25 24.63 ;
      RECT 31.07 21.69 31.23 24.63 ;
      RECT 33.59 21.69 33.75 24.63 ;
      RECT 31.07 21.69 33.75 21.85 ;
      RECT 32.67 36.47 34.55 36.63 ;
      RECT 34.39 35.86 34.55 36.63 ;
      RECT 33.53 35.23 33.69 36.63 ;
      RECT 32.67 35.86 32.83 36.63 ;
      RECT 34.49 35.23 34.65 36.05 ;
      RECT 32.57 35.23 32.73 36.05 ;
      RECT 34.49 37.11 34.65 38.19 ;
      RECT 33.53 36.79 33.69 38.19 ;
      RECT 32.57 37.11 32.73 38.19 ;
      RECT 34.39 36.79 34.55 37.39 ;
      RECT 32.67 36.79 32.83 37.39 ;
      RECT 32.67 36.79 34.55 36.95 ;
      RECT 34.45 21.37 34.61 23.37 ;
      RECT 30.61 21.37 34.61 21.53 ;
      RECT 33.96 20.73 34.12 21.53 ;
      RECT 30.61 20.78 30.77 21.53 ;
      RECT 33.29 50.66 33.45 51.5 ;
      RECT 33.29 50.66 34.09 50.82 ;
      RECT 33.93 50.18 34.09 50.82 ;
      RECT 33.93 50.18 34.57 50.5 ;
      RECT 34.41 47.07 34.57 50.5 ;
      RECT 34.09 47.07 34.57 47.23 ;
      RECT 34.09 45.44 34.25 47.23 ;
      RECT 34.41 56.67 34.57 61.86 ;
      RECT 33.13 56.67 34.57 56.83 ;
      RECT 34.25 54.4 34.41 56.83 ;
      RECT 33.13 56 33.29 56.83 ;
      RECT 34.09 47.39 34.25 49.72 ;
      RECT 33.77 47.39 34.25 47.55 ;
      RECT 33.77 43.85 33.93 47.55 ;
      RECT 33.77 43.85 34.55 44.01 ;
      RECT 34.39 39.56 34.55 44.01 ;
      RECT 34.21 39.56 34.55 39.84 ;
      RECT 34.21 39.16 34.37 39.84 ;
      RECT 32.99 53.23 33.27 53.51 ;
      RECT 33.11 53.03 33.27 53.51 ;
      RECT 33.11 53.03 34.09 53.19 ;
      RECT 33.93 50.98 34.09 53.19 ;
      RECT 33.93 52.54 34.13 52.82 ;
      RECT 33.93 50.98 34.47 51.14 ;
      RECT 34.25 50.8 34.47 51.14 ;
      RECT 32.65 68.07 34.47 68.23 ;
      RECT 34.31 62.02 34.47 68.23 ;
      RECT 34.09 62.02 34.47 62.18 ;
      RECT 34.09 57.45 34.25 62.18 ;
      RECT 32.65 57.45 34.25 57.61 ;
      RECT 32.65 57.39 32.97 57.61 ;
      RECT 32.81 53.74 32.97 57.61 ;
      RECT 32.65 51.32 32.81 53.9 ;
      RECT 32.65 51.32 33.13 51.48 ;
      RECT 32.97 49.88 33.13 51.48 ;
      RECT 32.97 49.88 33.45 50.04 ;
      RECT 33.29 47.71 33.45 50.04 ;
      RECT 33.29 47.71 33.91 47.99 ;
      RECT 33.93 54.06 34.09 56.51 ;
      RECT 33.93 54.06 34.45 54.22 ;
      RECT 34.29 51.34 34.45 54.22 ;
      RECT 34.25 52.98 34.45 54.22 ;
      RECT 34.25 51.34 34.45 52.12 ;
      RECT 33.14 18.78 34.26 18.94 ;
      RECT 34.08 17.48 34.26 18.94 ;
      RECT 32.18 17.26 32.35 18.8 ;
      RECT 32.19 16.12 32.35 18.8 ;
      RECT 31.22 16.44 31.38 18.8 ;
      RECT 33.14 16.03 33.3 18.94 ;
      RECT 31.17 16.44 31.38 17.57 ;
      RECT 34.08 16.44 34.24 18.94 ;
      RECT 31.17 17.26 32.35 17.42 ;
      RECT 31.17 16.44 31.45 17.42 ;
      RECT 33.95 14.52 34.11 16.71 ;
      RECT 30.17 16.12 33.3 16.28 ;
      RECT 32.99 14.52 33.15 16.28 ;
      RECT 31.99 14.84 32.15 16.28 ;
      RECT 32.99 14.52 34.11 14.68 ;
      RECT 33.89 34.44 34.23 34.72 ;
      RECT 33.89 32.44 34.05 34.72 ;
      RECT 33.89 33.11 34.23 33.39 ;
      RECT 33.89 32.44 34.23 32.72 ;
      RECT 33.89 40.7 34.23 40.98 ;
      RECT 33.89 38.7 34.05 40.98 ;
      RECT 33.89 40.03 34.23 40.31 ;
      RECT 33.89 38.7 34.23 38.98 ;
      RECT 34.05 21.85 34.21 24.3 ;
      RECT 33.91 21.85 34.21 22.13 ;
      RECT 33.89 24.79 34.09 25.35 ;
      RECT 33.89 24.79 34.21 25.03 ;
      RECT 32.57 28.04 32.89 28.32 ;
      RECT 32.73 25.99 32.89 28.32 ;
      RECT 33.92 27.02 34.08 27.7 ;
      RECT 32.73 27.02 34.08 27.18 ;
      RECT 32.73 25.99 33.11 26.23 ;
      RECT 32.95 25.16 33.11 26.23 ;
      RECT 32.59 20.26 32.75 21.05 ;
      RECT 32.59 20.26 33.32 20.44 ;
      RECT 33.16 19.89 33.32 20.44 ;
      RECT 33.16 19.89 33.98 20.05 ;
      RECT 33.79 19.61 33.98 20.05 ;
      RECT 33.79 19.61 34.07 19.77 ;
      RECT 33.53 55.68 33.69 56.51 ;
      RECT 33.29 55.68 33.69 55.84 ;
      RECT 33.29 53.67 33.45 55.84 ;
      RECT 33.29 53.67 33.93 53.83 ;
      RECT 33.65 53.35 33.93 53.83 ;
      RECT 33.39 51.7 33.77 51.92 ;
      RECT 33.61 50.98 33.77 51.92 ;
      RECT 32.97 52.58 33.73 52.86 ;
      RECT 33.57 52.18 33.73 52.86 ;
      RECT 32.97 51.64 33.13 52.86 ;
      RECT 33.27 12.53 33.43 13.61 ;
      RECT 33.43 11.88 33.59 12.69 ;
      RECT 32.47 11.77 32.71 12.05 ;
      RECT 32.47 11.88 33.59 12.04 ;
      RECT 33.35 8.88 33.51 12.04 ;
      RECT 33.29 62.9 33.45 67.89 ;
      RECT 33.29 65.82 33.51 66.55 ;
      RECT 32.97 47.39 33.13 49.72 ;
      RECT 32.97 47.39 33.45 47.55 ;
      RECT 33.29 43.85 33.45 47.55 ;
      RECT 32.67 43.85 33.45 44.01 ;
      RECT 32.67 39.56 32.83 44.01 ;
      RECT 32.67 39.56 33.01 39.84 ;
      RECT 32.85 39.16 33.01 39.84 ;
      RECT 33.27 22.01 33.43 23.37 ;
      RECT 32.65 22.01 33.43 22.17 ;
      RECT 32.95 24.72 33.33 24.96 ;
      RECT 32.95 22.35 33.11 24.96 ;
      RECT 32.99 34.44 33.33 34.72 ;
      RECT 33.17 32.44 33.33 34.72 ;
      RECT 32.99 33.11 33.33 33.39 ;
      RECT 32.99 32.44 33.33 32.72 ;
      RECT 32.99 40.7 33.33 40.98 ;
      RECT 33.17 38.7 33.33 40.98 ;
      RECT 32.99 40.03 33.33 40.31 ;
      RECT 32.99 38.7 33.33 38.98 ;
      RECT 31.69 12.21 31.85 13.28 ;
      RECT 31.69 12.21 33.27 12.37 ;
      RECT 32.15 11.47 32.31 12.37 ;
      RECT 32.21 10.85 32.37 11.63 ;
      RECT 32.81 62.9 32.97 67.89 ;
      RECT 32.81 64.59 33.09 65.31 ;
      RECT 32.33 46.75 32.49 47.43 ;
      RECT 32.01 46.75 32.81 46.91 ;
      RECT 32.65 44.23 32.81 46.91 ;
      RECT 32.01 44.23 32.17 46.91 ;
      RECT 32.53 10.51 32.69 11.24 ;
      RECT 32.03 10.51 32.69 10.67 ;
      RECT 32.38 8.96 32.54 9.79 ;
      RECT 31.35 8.96 32.54 9.12 ;
      RECT 32.05 20.63 32.33 20.79 ;
      RECT 32.17 19.59 32.33 20.79 ;
      RECT 30.11 34.88 32.31 35.04 ;
      RECT 32.03 34.59 32.31 35.04 ;
      RECT 31.09 34.59 31.33 35.04 ;
      RECT 30.11 34.59 30.39 35.04 ;
      RECT 31.09 38.38 31.33 39.02 ;
      RECT 32.03 38.38 32.31 38.83 ;
      RECT 30.11 38.38 30.39 38.83 ;
      RECT 30.11 38.38 32.31 38.54 ;
      RECT 31.93 28.04 32.25 28.32 ;
      RECT 31.93 25.99 32.09 28.32 ;
      RECT 30.74 27.02 30.9 27.7 ;
      RECT 30.74 27.02 32.09 27.18 ;
      RECT 31.71 25.99 32.09 26.23 ;
      RECT 31.71 25.16 31.87 26.23 ;
      RECT 30.27 36.47 32.15 36.63 ;
      RECT 31.99 35.88 32.15 36.63 ;
      RECT 31.13 35.23 31.29 36.63 ;
      RECT 30.27 35.88 30.43 36.63 ;
      RECT 32.09 35.23 32.25 36.06 ;
      RECT 30.17 35.23 30.33 36.06 ;
      RECT 32.09 37.11 32.25 38.19 ;
      RECT 31.13 36.79 31.29 38.19 ;
      RECT 30.17 37.11 30.33 38.19 ;
      RECT 31.99 36.79 32.15 37.39 ;
      RECT 30.27 36.79 30.43 37.39 ;
      RECT 30.27 36.79 32.15 36.95 ;
      RECT 31.39 22.01 31.55 23.37 ;
      RECT 31.39 22.01 32.17 22.17 ;
      RECT 30.35 68.07 32.17 68.23 ;
      RECT 30.35 62.02 30.51 68.23 ;
      RECT 30.35 62.02 30.73 62.18 ;
      RECT 30.57 57.45 30.73 62.18 ;
      RECT 30.57 57.45 32.17 57.61 ;
      RECT 31.85 57.39 32.17 57.61 ;
      RECT 31.85 53.74 32.01 57.61 ;
      RECT 32.01 51.32 32.17 53.9 ;
      RECT 31.69 51.32 32.17 51.48 ;
      RECT 31.69 49.88 31.85 51.48 ;
      RECT 31.37 49.88 31.85 50.04 ;
      RECT 31.37 47.71 31.53 50.04 ;
      RECT 30.91 47.71 31.53 47.99 ;
      RECT 31.69 47.39 31.85 49.72 ;
      RECT 31.37 47.39 31.85 47.55 ;
      RECT 31.37 43.85 31.53 47.55 ;
      RECT 31.37 43.85 32.15 44.01 ;
      RECT 31.99 39.56 32.15 44.01 ;
      RECT 31.81 39.56 32.15 39.84 ;
      RECT 31.81 39.16 31.97 39.84 ;
      RECT 31.51 14.44 31.67 15.64 ;
      RECT 31.51 14.44 32.01 14.6 ;
      RECT 31.85 62.9 32.01 67.89 ;
      RECT 31.73 64.59 32.01 65.31 ;
      RECT 31.49 24.72 31.87 24.96 ;
      RECT 31.71 22.35 31.87 24.96 ;
      RECT 31.21 12.32 31.37 13.37 ;
      RECT 31.33 11.56 31.49 12.48 ;
      RECT 30.73 11.56 31.85 11.72 ;
      RECT 31.69 10.27 31.85 11.72 ;
      RECT 30.73 10.4 30.89 11.72 ;
      RECT 31.09 52.58 31.85 52.86 ;
      RECT 31.69 51.64 31.85 52.86 ;
      RECT 31.09 52.18 31.25 52.86 ;
      RECT 31.49 34.44 31.83 34.72 ;
      RECT 31.49 32.44 31.65 34.72 ;
      RECT 31.49 33.11 31.83 33.39 ;
      RECT 31.49 32.44 31.83 32.72 ;
      RECT 31.49 40.7 31.83 40.98 ;
      RECT 31.49 38.7 31.65 40.98 ;
      RECT 31.49 40.03 31.83 40.31 ;
      RECT 31.49 38.7 31.83 38.98 ;
      RECT 31.55 53.23 31.83 53.51 ;
      RECT 31.55 53.03 31.71 53.51 ;
      RECT 30.73 53.03 31.71 53.19 ;
      RECT 30.73 50.98 30.89 53.19 ;
      RECT 30.69 52.54 30.89 52.82 ;
      RECT 30.35 50.98 30.89 51.14 ;
      RECT 30.35 50.8 30.57 51.14 ;
      RECT 30.25 56.67 30.41 61.86 ;
      RECT 30.25 56.67 31.69 56.83 ;
      RECT 31.53 56 31.69 56.83 ;
      RECT 30.41 54.4 30.57 56.83 ;
      RECT 31.39 26.36 31.55 26.72 ;
      RECT 29.25 26.36 31.55 26.52 ;
      RECT 29.25 26.04 29.41 26.52 ;
      RECT 28.6 26.04 29.41 26.2 ;
      RECT 31.37 50.66 31.53 51.5 ;
      RECT 30.73 50.66 31.53 50.82 ;
      RECT 30.73 50.18 30.89 50.82 ;
      RECT 30.25 50.18 30.89 50.5 ;
      RECT 30.25 47.07 30.41 50.5 ;
      RECT 30.25 47.07 30.73 47.23 ;
      RECT 30.57 45.44 30.73 47.23 ;
      RECT 31.13 55.68 31.29 56.51 ;
      RECT 31.13 55.68 31.53 55.84 ;
      RECT 31.37 53.67 31.53 55.84 ;
      RECT 30.89 53.67 31.53 53.83 ;
      RECT 30.89 53.35 31.17 53.83 ;
      RECT 31.37 62.9 31.53 67.89 ;
      RECT 31.31 65.82 31.53 66.55 ;
      RECT 31.05 51.7 31.43 51.92 ;
      RECT 31.05 50.98 31.21 51.92 ;
      RECT 29.22 28.01 31.38 28.17 ;
      RECT 31.22 27.34 31.38 28.17 ;
      RECT 31.06 27.93 31.38 28.17 ;
      RECT 30.22 26.97 30.38 28.17 ;
      RECT 29.22 26.68 29.38 28.17 ;
      RECT 30.73 12 30.89 12.84 ;
      RECT 30.73 12 31.17 12.16 ;
      RECT 31.01 11.88 31.17 12.16 ;
      RECT 29.48 8.82 31.07 8.98 ;
      RECT 30.91 7.16 31.07 8.98 ;
      RECT 30.57 47.39 30.73 49.72 ;
      RECT 30.57 47.39 31.05 47.55 ;
      RECT 30.89 43.85 31.05 47.55 ;
      RECT 30.27 43.85 31.05 44.01 ;
      RECT 30.27 39.56 30.43 44.01 ;
      RECT 30.27 39.56 30.61 39.84 ;
      RECT 30.45 39.16 30.61 39.84 ;
      RECT 30.88 9.92 31.04 10.24 ;
      RECT 30.64 9.92 31.04 10.12 ;
      RECT 29.85 15.8 30.01 17.77 ;
      RECT 29.85 15.8 30.67 15.96 ;
      RECT 30.67 14.42 30.83 15.88 ;
      RECT 30.49 15.72 30.83 15.88 ;
      RECT 30.67 14.42 31.01 14.58 ;
      RECT 30.73 24.79 30.93 25.35 ;
      RECT 30.61 24.79 30.93 25.03 ;
      RECT 30.59 34.44 30.93 34.72 ;
      RECT 30.77 32.44 30.93 34.72 ;
      RECT 30.59 33.11 30.93 33.39 ;
      RECT 30.59 32.44 30.93 32.72 ;
      RECT 30.59 40.7 30.93 40.98 ;
      RECT 30.77 38.7 30.93 40.98 ;
      RECT 30.59 40.03 30.93 40.31 ;
      RECT 30.59 38.7 30.93 38.98 ;
      RECT 30.61 21.85 30.77 24.3 ;
      RECT 30.61 21.85 30.91 22.13 ;
      RECT 30.73 54.06 30.89 56.51 ;
      RECT 30.37 54.06 30.89 54.22 ;
      RECT 30.37 52.98 30.57 54.22 ;
      RECT 30.37 51.34 30.53 54.22 ;
      RECT 30.37 51.34 30.57 52.12 ;
      RECT 30.23 18.51 30.42 18.94 ;
      RECT 30.03 18.51 30.72 18.7 ;
      RECT 30.21 21.29 30.37 23.37 ;
      RECT 30.29 19.81 30.45 21.46 ;
      RECT 29.83 12.58 30.11 13.24 ;
      RECT 29.95 11.84 30.11 13.24 ;
      RECT 29.59 11.84 29.75 12.12 ;
      RECT 29.59 11.84 30.43 12 ;
      RECT 30.27 10.46 30.43 12 ;
      RECT 29.93 46.75 30.09 47.43 ;
      RECT 29.61 46.75 30.41 46.91 ;
      RECT 30.25 44.23 30.41 46.91 ;
      RECT 29.61 44.23 29.77 46.91 ;
      RECT 29.77 26.02 30.33 26.18 ;
      RECT 29.77 25.58 29.93 26.18 ;
      RECT 29.23 25.58 29.93 25.74 ;
      RECT 29.23 24 29.43 25.74 ;
      RECT 28.49 24.24 29.43 24.52 ;
      RECT 28.49 21.85 28.65 24.52 ;
      RECT 29.16 9.14 29.35 9.52 ;
      RECT 29.16 9.14 30.29 9.3 ;
      RECT 29.16 8.52 29.32 9.52 ;
      RECT 29.14 8.36 29.3 8.64 ;
      RECT 29.53 18.13 30.19 18.3 ;
      RECT 29.53 15 29.69 18.3 ;
      RECT 29.53 15.32 30.23 15.64 ;
      RECT 29.07 15 29.69 15.16 ;
      RECT 29.79 9.68 29.95 11.68 ;
      RECT 25.27 9.68 25.43 11.68 ;
      RECT 28.33 9.68 28.49 11.36 ;
      RECT 26.73 9.68 26.89 11.36 ;
      RECT 26.73 10.76 28.49 10.92 ;
      RECT 27.53 8.38 27.69 10.92 ;
      RECT 28.33 9.68 29.95 9.84 ;
      RECT 29.67 9.46 29.83 9.84 ;
      RECT 25.27 9.68 26.89 9.84 ;
      RECT 25.39 9.46 25.55 9.84 ;
      RECT 29.74 26.68 29.9 27.85 ;
      RECT 29.7 26.68 29.94 27.33 ;
      RECT 27.71 34.88 29.91 35.04 ;
      RECT 29.63 34.59 29.91 35.04 ;
      RECT 28.69 34.59 28.93 35.04 ;
      RECT 27.71 34.59 27.99 35.04 ;
      RECT 28.69 38.38 28.93 39.02 ;
      RECT 29.63 38.38 29.91 38.83 ;
      RECT 27.71 38.38 27.99 38.83 ;
      RECT 27.71 38.38 29.91 38.54 ;
      RECT 29.69 13.5 29.85 14.2 ;
      RECT 29.51 13.5 29.85 13.66 ;
      RECT 29.51 12.52 29.67 13.66 ;
      RECT 29.27 12.52 29.67 12.84 ;
      RECT 29.27 10.84 29.43 12.84 ;
      RECT 27.87 36.47 29.75 36.63 ;
      RECT 29.59 35.86 29.75 36.63 ;
      RECT 28.73 35.23 28.89 36.63 ;
      RECT 27.87 35.86 28.03 36.63 ;
      RECT 29.69 35.23 29.85 36.05 ;
      RECT 27.77 35.23 27.93 36.05 ;
      RECT 29.69 37.11 29.85 38.19 ;
      RECT 28.73 36.79 28.89 38.19 ;
      RECT 27.77 37.11 27.93 38.19 ;
      RECT 29.59 36.79 29.75 37.39 ;
      RECT 27.87 36.79 28.03 37.39 ;
      RECT 27.87 36.79 29.75 36.95 ;
      RECT 28.49 50.66 28.65 51.5 ;
      RECT 28.49 50.66 29.29 50.82 ;
      RECT 29.13 50.18 29.29 50.82 ;
      RECT 29.13 50.18 29.77 50.5 ;
      RECT 29.61 47.07 29.77 50.5 ;
      RECT 29.29 47.07 29.77 47.23 ;
      RECT 29.29 45.44 29.45 47.23 ;
      RECT 29.61 56.67 29.77 61.86 ;
      RECT 28.33 56.67 29.77 56.83 ;
      RECT 29.45 54.4 29.61 56.83 ;
      RECT 28.33 56 28.49 56.83 ;
      RECT 29.29 47.39 29.45 49.72 ;
      RECT 28.97 47.39 29.45 47.55 ;
      RECT 28.97 43.85 29.13 47.55 ;
      RECT 28.97 43.85 29.75 44.01 ;
      RECT 29.59 39.56 29.75 44.01 ;
      RECT 29.41 39.56 29.75 39.84 ;
      RECT 29.41 39.16 29.57 39.84 ;
      RECT 29.55 23.12 29.71 23.84 ;
      RECT 28.81 23.12 29.71 23.28 ;
      RECT 28.81 20.86 28.97 23.28 ;
      RECT 28.81 20.86 29.17 21.02 ;
      RECT 29.01 20.74 29.17 21.02 ;
      RECT 28.2 28.52 29.29 28.68 ;
      RECT 29.01 28.35 29.29 28.68 ;
      RECT 29.01 28.35 29.69 28.51 ;
      RECT 28.19 53.23 28.47 53.51 ;
      RECT 28.31 53.03 28.47 53.51 ;
      RECT 28.31 53.03 29.29 53.19 ;
      RECT 29.13 50.98 29.29 53.19 ;
      RECT 29.13 52.54 29.33 52.82 ;
      RECT 29.13 50.98 29.67 51.14 ;
      RECT 29.45 50.8 29.67 51.14 ;
      RECT 27.85 68.07 29.67 68.23 ;
      RECT 29.51 62.02 29.67 68.23 ;
      RECT 29.29 62.02 29.67 62.18 ;
      RECT 29.29 57.45 29.45 62.18 ;
      RECT 27.85 57.45 29.45 57.61 ;
      RECT 27.85 57.39 28.17 57.61 ;
      RECT 28.01 53.74 28.17 57.61 ;
      RECT 27.85 51.32 28.01 53.9 ;
      RECT 27.85 51.32 28.33 51.48 ;
      RECT 28.17 49.88 28.33 51.48 ;
      RECT 28.17 49.88 28.65 50.04 ;
      RECT 28.49 47.71 28.65 50.04 ;
      RECT 28.49 47.71 29.11 47.99 ;
      RECT 29.13 54.06 29.29 56.51 ;
      RECT 29.13 54.06 29.65 54.22 ;
      RECT 29.49 51.34 29.65 54.22 ;
      RECT 29.45 52.98 29.65 54.22 ;
      RECT 29.45 51.34 29.65 52.12 ;
      RECT 29.09 13.06 29.25 13.54 ;
      RECT 28.81 13.06 29.25 13.22 ;
      RECT 28.81 10 28.97 13.22 ;
      RECT 28.81 10 29.63 10.16 ;
      RECT 29.17 22.29 29.41 22.53 ;
      RECT 29.17 21.18 29.33 22.53 ;
      RECT 29.13 21.18 29.33 21.58 ;
      RECT 29.33 19.81 29.5 21.35 ;
      RECT 29.09 34.44 29.43 34.72 ;
      RECT 29.09 32.44 29.25 34.72 ;
      RECT 29.09 33.11 29.43 33.39 ;
      RECT 29.09 32.44 29.43 32.72 ;
      RECT 29.09 40.7 29.43 40.98 ;
      RECT 29.09 38.7 29.25 40.98 ;
      RECT 29.09 40.03 29.43 40.31 ;
      RECT 29.09 38.7 29.43 38.98 ;
      RECT 28.97 17.24 29.13 19 ;
      RECT 28.01 14.39 28.17 18.85 ;
      RECT 28.01 17.24 29.13 17.4 ;
      RECT 27.99 15.32 28.19 16.04 ;
      RECT 28.01 14.39 28.19 16.04 ;
      RECT 28.73 55.68 28.89 56.51 ;
      RECT 28.49 55.68 28.89 55.84 ;
      RECT 28.49 53.67 28.65 55.84 ;
      RECT 28.49 53.67 29.13 53.83 ;
      RECT 28.85 53.35 29.13 53.83 ;
      RECT 28.28 24.7 28.44 28.32 ;
      RECT 28.28 25.16 28.97 25.32 ;
      RECT 27.75 24.7 28.44 24.86 ;
      RECT 28.59 51.7 28.97 51.92 ;
      RECT 28.81 50.98 28.97 51.92 ;
      RECT 28.17 52.58 28.93 52.86 ;
      RECT 28.77 52.18 28.93 52.86 ;
      RECT 28.17 51.64 28.33 52.86 ;
      RECT 28.49 62.9 28.65 67.89 ;
      RECT 28.49 65.82 28.71 66.55 ;
      RECT 27.93 9.36 28.09 10.6 ;
      RECT 27.93 9.36 28.67 9.52 ;
      RECT 28.17 47.39 28.33 49.72 ;
      RECT 28.17 47.39 28.65 47.55 ;
      RECT 28.49 43.85 28.65 47.55 ;
      RECT 27.87 43.85 28.65 44.01 ;
      RECT 27.87 39.56 28.03 44.01 ;
      RECT 27.87 39.56 28.21 39.84 ;
      RECT 28.05 39.16 28.21 39.84 ;
      RECT 28.19 34.44 28.53 34.72 ;
      RECT 28.37 32.44 28.53 34.72 ;
      RECT 28.19 33.11 28.53 33.39 ;
      RECT 28.19 32.44 28.53 32.72 ;
      RECT 28.19 40.7 28.53 40.98 ;
      RECT 28.37 38.7 28.53 40.98 ;
      RECT 28.19 40.03 28.53 40.31 ;
      RECT 28.19 38.7 28.53 38.98 ;
      RECT 28.09 11.52 28.25 12.43 ;
      RECT 28.09 11.75 28.33 12.03 ;
      RECT 27.81 11.52 28.25 11.68 ;
      RECT 27.81 11.08 27.97 11.68 ;
      RECT 28.01 62.9 28.17 67.89 ;
      RECT 28.01 64.59 28.29 65.31 ;
      RECT 28.01 23.73 28.19 24.54 ;
      RECT 28.01 20.48 28.17 24.54 ;
      RECT 27.53 46.75 27.69 47.43 ;
      RECT 27.21 46.75 28.01 46.91 ;
      RECT 27.85 44.23 28.01 46.91 ;
      RECT 27.21 44.23 27.37 46.91 ;
      RECT 27.8 26.15 27.96 28.96 ;
      RECT 27.77 26.15 27.96 26.51 ;
      RECT 25.31 34.88 27.51 35.04 ;
      RECT 27.23 34.59 27.51 35.04 ;
      RECT 26.29 34.59 26.53 35.04 ;
      RECT 25.31 34.59 25.59 35.04 ;
      RECT 26.29 38.38 26.53 39.02 ;
      RECT 27.23 38.38 27.51 38.83 ;
      RECT 25.31 38.38 25.59 38.83 ;
      RECT 25.31 38.38 27.51 38.54 ;
      RECT 26.78 24.7 26.94 28.32 ;
      RECT 26.25 25.16 26.94 25.32 ;
      RECT 26.78 24.7 27.47 24.86 ;
      RECT 27.26 26.15 27.42 28.96 ;
      RECT 27.26 26.15 27.45 26.51 ;
      RECT 25.47 36.47 27.35 36.63 ;
      RECT 27.19 35.88 27.35 36.63 ;
      RECT 26.33 35.23 26.49 36.63 ;
      RECT 25.47 35.88 25.63 36.63 ;
      RECT 27.29 35.23 27.45 36.06 ;
      RECT 25.37 35.23 25.53 36.06 ;
      RECT 27.29 37.11 27.45 38.19 ;
      RECT 26.33 36.79 26.49 38.19 ;
      RECT 25.37 37.11 25.53 38.19 ;
      RECT 27.19 36.79 27.35 37.39 ;
      RECT 25.47 36.79 25.63 37.39 ;
      RECT 25.47 36.79 27.35 36.95 ;
      RECT 26.97 11.52 27.13 12.43 ;
      RECT 26.89 11.75 27.13 12.03 ;
      RECT 26.97 11.52 27.41 11.68 ;
      RECT 27.25 11.08 27.41 11.68 ;
      RECT 25.55 68.07 27.37 68.23 ;
      RECT 25.55 62.02 25.71 68.23 ;
      RECT 25.55 62.02 25.93 62.18 ;
      RECT 25.77 57.45 25.93 62.18 ;
      RECT 25.77 57.45 27.37 57.61 ;
      RECT 27.05 57.39 27.37 57.61 ;
      RECT 27.05 53.74 27.21 57.61 ;
      RECT 27.21 51.32 27.37 53.9 ;
      RECT 26.89 51.32 27.37 51.48 ;
      RECT 26.89 49.88 27.05 51.48 ;
      RECT 26.57 49.88 27.05 50.04 ;
      RECT 26.57 47.71 26.73 50.04 ;
      RECT 26.11 47.71 26.73 47.99 ;
      RECT 26.89 47.39 27.05 49.72 ;
      RECT 26.57 47.39 27.05 47.55 ;
      RECT 26.57 43.85 26.73 47.55 ;
      RECT 26.57 43.85 27.35 44.01 ;
      RECT 27.19 39.56 27.35 44.01 ;
      RECT 27.01 39.56 27.35 39.84 ;
      RECT 27.01 39.16 27.17 39.84 ;
      RECT 27.13 9.36 27.29 10.6 ;
      RECT 26.55 9.36 27.29 9.52 ;
      RECT 26.09 17.24 26.25 19 ;
      RECT 27.05 14.39 27.21 18.85 ;
      RECT 26.09 17.24 27.21 17.4 ;
      RECT 27.03 15.32 27.23 16.04 ;
      RECT 27.03 14.39 27.21 16.04 ;
      RECT 27.03 23.73 27.21 24.54 ;
      RECT 27.05 20.48 27.21 24.54 ;
      RECT 27.05 62.9 27.21 67.89 ;
      RECT 26.93 64.59 27.21 65.31 ;
      RECT 26.29 52.58 27.05 52.86 ;
      RECT 26.89 51.64 27.05 52.86 ;
      RECT 26.29 52.18 26.45 52.86 ;
      RECT 26.69 34.44 27.03 34.72 ;
      RECT 26.69 32.44 26.85 34.72 ;
      RECT 26.69 33.11 27.03 33.39 ;
      RECT 26.69 32.44 27.03 32.72 ;
      RECT 26.69 40.7 27.03 40.98 ;
      RECT 26.69 38.7 26.85 40.98 ;
      RECT 26.69 40.03 27.03 40.31 ;
      RECT 26.69 38.7 27.03 38.98 ;
      RECT 26.75 53.23 27.03 53.51 ;
      RECT 26.75 53.03 26.91 53.51 ;
      RECT 25.93 53.03 26.91 53.19 ;
      RECT 25.93 50.98 26.09 53.19 ;
      RECT 25.89 52.54 26.09 52.82 ;
      RECT 25.55 50.98 26.09 51.14 ;
      RECT 25.55 50.8 25.77 51.14 ;
      RECT 25.93 28.52 27.02 28.68 ;
      RECT 25.93 28.35 26.21 28.68 ;
      RECT 25.53 28.35 26.21 28.51 ;
      RECT 25.45 56.67 25.61 61.86 ;
      RECT 25.45 56.67 26.89 56.83 ;
      RECT 26.73 56 26.89 56.83 ;
      RECT 25.61 54.4 25.77 56.83 ;
      RECT 24.89 26.02 25.45 26.18 ;
      RECT 25.29 25.58 25.45 26.18 ;
      RECT 25.29 25.58 25.99 25.74 ;
      RECT 25.79 24 25.99 25.74 ;
      RECT 25.79 24.24 26.73 24.52 ;
      RECT 26.57 21.85 26.73 24.52 ;
      RECT 26.57 50.66 26.73 51.5 ;
      RECT 25.93 50.66 26.73 50.82 ;
      RECT 25.93 50.18 26.09 50.82 ;
      RECT 25.45 50.18 26.09 50.5 ;
      RECT 25.45 47.07 25.61 50.5 ;
      RECT 25.45 47.07 25.93 47.23 ;
      RECT 25.77 45.44 25.93 47.23 ;
      RECT 26.33 55.68 26.49 56.51 ;
      RECT 26.33 55.68 26.73 55.84 ;
      RECT 26.57 53.67 26.73 55.84 ;
      RECT 26.09 53.67 26.73 53.83 ;
      RECT 26.09 53.35 26.37 53.83 ;
      RECT 26.57 62.9 26.73 67.89 ;
      RECT 26.51 65.82 26.73 66.55 ;
      RECT 26.25 51.7 26.63 51.92 ;
      RECT 26.25 50.98 26.41 51.92 ;
      RECT 23.67 26.36 23.83 26.72 ;
      RECT 23.67 26.36 25.97 26.52 ;
      RECT 25.81 26.04 25.97 26.52 ;
      RECT 25.81 26.04 26.62 26.2 ;
      RECT 25.97 13.06 26.13 13.54 ;
      RECT 25.97 13.06 26.41 13.22 ;
      RECT 26.25 10 26.41 13.22 ;
      RECT 25.59 10 26.41 10.16 ;
      RECT 25.51 23.12 25.67 23.84 ;
      RECT 25.51 23.12 26.41 23.28 ;
      RECT 26.25 20.86 26.41 23.28 ;
      RECT 26.05 20.86 26.41 21.02 ;
      RECT 26.05 20.74 26.21 21.02 ;
      RECT 25.77 47.39 25.93 49.72 ;
      RECT 25.77 47.39 26.25 47.55 ;
      RECT 26.09 43.85 26.25 47.55 ;
      RECT 25.47 43.85 26.25 44.01 ;
      RECT 25.47 39.56 25.63 44.01 ;
      RECT 25.47 39.56 25.81 39.84 ;
      RECT 25.65 39.16 25.81 39.84 ;
      RECT 25.03 18.13 25.69 18.3 ;
      RECT 25.53 15 25.69 18.3 ;
      RECT 24.99 15.32 25.69 15.64 ;
      RECT 25.53 15 26.15 15.16 ;
      RECT 25.79 34.44 26.13 34.72 ;
      RECT 25.97 32.44 26.13 34.72 ;
      RECT 25.79 33.11 26.13 33.39 ;
      RECT 25.79 32.44 26.13 32.72 ;
      RECT 25.79 40.7 26.13 40.98 ;
      RECT 25.97 38.7 26.13 40.98 ;
      RECT 25.79 40.03 26.13 40.31 ;
      RECT 25.79 38.7 26.13 38.98 ;
      RECT 25.81 22.29 26.05 22.53 ;
      RECT 25.89 21.18 26.05 22.53 ;
      RECT 25.89 21.18 26.09 21.58 ;
      RECT 25.72 19.81 25.89 21.35 ;
      RECT 25.93 54.06 26.09 56.51 ;
      RECT 25.57 54.06 26.09 54.22 ;
      RECT 25.57 52.98 25.77 54.22 ;
      RECT 25.57 51.34 25.73 54.22 ;
      RECT 25.57 51.34 25.77 52.12 ;
      RECT 25.87 9.14 26.06 9.52 ;
      RECT 24.93 9.14 26.06 9.3 ;
      RECT 25.9 8.52 26.06 9.52 ;
      RECT 25.92 8.36 26.08 8.64 ;
      RECT 23.84 28.01 26 28.17 ;
      RECT 25.84 26.68 26 28.17 ;
      RECT 24.84 26.97 25 28.17 ;
      RECT 23.84 27.93 24.16 28.17 ;
      RECT 23.84 27.34 24 28.17 ;
      RECT 25.37 13.5 25.53 14.2 ;
      RECT 25.37 13.5 25.71 13.66 ;
      RECT 25.55 12.52 25.71 13.66 ;
      RECT 25.55 12.52 25.95 12.84 ;
      RECT 25.79 10.84 25.95 12.84 ;
      RECT 24.15 8.82 25.74 8.98 ;
      RECT 24.15 7.16 24.31 8.98 ;
      RECT 25.11 12.58 25.39 13.24 ;
      RECT 25.11 11.84 25.27 13.24 ;
      RECT 25.47 11.84 25.63 12.12 ;
      RECT 24.79 11.84 25.63 12 ;
      RECT 24.79 10.46 24.95 12 ;
      RECT 25.13 46.75 25.29 47.43 ;
      RECT 24.81 46.75 25.61 46.91 ;
      RECT 25.45 44.23 25.61 46.91 ;
      RECT 24.81 44.23 24.97 46.91 ;
      RECT 25.32 26.68 25.48 27.85 ;
      RECT 25.28 26.68 25.52 27.33 ;
      RECT 25.21 15.8 25.37 17.77 ;
      RECT 24.55 15.8 25.37 15.96 ;
      RECT 24.39 14.42 24.55 15.88 ;
      RECT 24.39 15.72 24.73 15.88 ;
      RECT 24.21 14.42 24.55 14.58 ;
      RECT 20.25 28.74 25.37 28.9 ;
      RECT 23.45 27.92 23.61 28.9 ;
      RECT 22.01 27.92 22.17 28.9 ;
      RECT 24.8 18.51 24.99 18.94 ;
      RECT 24.5 18.51 25.19 18.7 ;
      RECT 22.91 34.88 25.11 35.04 ;
      RECT 24.83 34.59 25.11 35.04 ;
      RECT 23.89 34.59 24.13 35.04 ;
      RECT 22.91 34.59 23.19 35.04 ;
      RECT 23.89 38.38 24.13 39.02 ;
      RECT 24.83 38.38 25.11 38.83 ;
      RECT 22.91 38.38 23.19 38.83 ;
      RECT 22.91 38.38 25.11 38.54 ;
      RECT 22.73 21.69 22.89 26.21 ;
      RECT 23.97 24.35 24.13 26.2 ;
      RECT 21.49 24.34 21.65 26.2 ;
      RECT 24.85 24.04 25.07 25.52 ;
      RECT 20.55 24.04 20.77 25.52 ;
      RECT 23.97 24.46 25.07 24.63 ;
      RECT 20.55 24.46 21.65 24.63 ;
      RECT 21.47 21.69 21.63 24.63 ;
      RECT 23.99 21.69 24.15 24.63 ;
      RECT 21.47 21.69 24.15 21.85 ;
      RECT 20.96 18.78 22.08 18.94 ;
      RECT 23.84 16.44 24 18.8 ;
      RECT 22.87 17.26 23.04 18.8 ;
      RECT 21.92 16.03 22.08 18.94 ;
      RECT 20.96 17.48 21.14 18.94 ;
      RECT 23.84 16.44 24.05 17.57 ;
      RECT 20.98 16.44 21.14 18.94 ;
      RECT 22.87 17.26 24.05 17.42 ;
      RECT 23.77 16.44 24.05 17.42 ;
      RECT 22.87 16.12 23.03 18.8 ;
      RECT 21.11 14.52 21.27 16.71 ;
      RECT 21.92 16.12 25.05 16.28 ;
      RECT 23.07 14.84 23.23 16.28 ;
      RECT 22.07 14.52 22.23 16.28 ;
      RECT 21.11 14.52 22.23 14.68 ;
      RECT 23.07 36.47 24.95 36.63 ;
      RECT 24.79 35.86 24.95 36.63 ;
      RECT 23.93 35.23 24.09 36.63 ;
      RECT 23.07 35.86 23.23 36.63 ;
      RECT 24.89 35.23 25.05 36.05 ;
      RECT 22.97 35.23 23.13 36.05 ;
      RECT 24.89 37.11 25.05 38.19 ;
      RECT 23.93 36.79 24.09 38.19 ;
      RECT 22.97 37.11 23.13 38.19 ;
      RECT 24.79 36.79 24.95 37.39 ;
      RECT 23.07 36.79 23.23 37.39 ;
      RECT 23.07 36.79 24.95 36.95 ;
      RECT 24.85 21.29 25.01 23.37 ;
      RECT 24.77 19.81 24.93 21.46 ;
      RECT 23.69 50.66 23.85 51.5 ;
      RECT 23.69 50.66 24.49 50.82 ;
      RECT 24.33 50.18 24.49 50.82 ;
      RECT 24.33 50.18 24.97 50.5 ;
      RECT 24.81 47.07 24.97 50.5 ;
      RECT 24.49 47.07 24.97 47.23 ;
      RECT 24.49 45.44 24.65 47.23 ;
      RECT 24.81 56.67 24.97 61.86 ;
      RECT 23.53 56.67 24.97 56.83 ;
      RECT 24.65 54.4 24.81 56.83 ;
      RECT 23.53 56 23.69 56.83 ;
      RECT 24.49 47.39 24.65 49.72 ;
      RECT 24.17 47.39 24.65 47.55 ;
      RECT 24.17 43.85 24.33 47.55 ;
      RECT 24.17 43.85 24.95 44.01 ;
      RECT 24.79 39.56 24.95 44.01 ;
      RECT 24.61 39.56 24.95 39.84 ;
      RECT 24.61 39.16 24.77 39.84 ;
      RECT 23.39 53.23 23.67 53.51 ;
      RECT 23.51 53.03 23.67 53.51 ;
      RECT 23.51 53.03 24.49 53.19 ;
      RECT 24.33 50.98 24.49 53.19 ;
      RECT 24.33 52.54 24.53 52.82 ;
      RECT 24.33 50.98 24.87 51.14 ;
      RECT 24.65 50.8 24.87 51.14 ;
      RECT 23.05 68.07 24.87 68.23 ;
      RECT 24.71 62.02 24.87 68.23 ;
      RECT 24.49 62.02 24.87 62.18 ;
      RECT 24.49 57.45 24.65 62.18 ;
      RECT 23.05 57.45 24.65 57.61 ;
      RECT 23.05 57.39 23.37 57.61 ;
      RECT 23.21 53.74 23.37 57.61 ;
      RECT 23.05 51.32 23.21 53.9 ;
      RECT 23.05 51.32 23.53 51.48 ;
      RECT 23.37 49.88 23.53 51.48 ;
      RECT 23.37 49.88 23.85 50.04 ;
      RECT 23.69 47.71 23.85 50.04 ;
      RECT 23.69 47.71 24.31 47.99 ;
      RECT 24.33 54.06 24.49 56.51 ;
      RECT 24.33 54.06 24.85 54.22 ;
      RECT 24.69 51.34 24.85 54.22 ;
      RECT 24.65 52.98 24.85 54.22 ;
      RECT 24.65 51.34 24.85 52.12 ;
      RECT 24.29 34.44 24.63 34.72 ;
      RECT 24.29 32.44 24.45 34.72 ;
      RECT 24.29 33.11 24.63 33.39 ;
      RECT 24.29 32.44 24.63 32.72 ;
      RECT 24.29 40.7 24.63 40.98 ;
      RECT 24.29 38.7 24.45 40.98 ;
      RECT 24.29 40.03 24.63 40.31 ;
      RECT 24.29 38.7 24.63 38.98 ;
      RECT 20.61 21.37 20.77 23.37 ;
      RECT 20.61 21.37 24.61 21.53 ;
      RECT 24.45 20.78 24.61 21.53 ;
      RECT 21.1 20.73 21.26 21.53 ;
      RECT 24.45 21.85 24.61 24.3 ;
      RECT 24.31 21.85 24.61 22.13 ;
      RECT 24.29 24.79 24.49 25.35 ;
      RECT 24.29 24.79 24.61 25.03 ;
      RECT 24.18 9.92 24.34 10.24 ;
      RECT 24.18 9.92 24.58 10.12 ;
      RECT 23.85 12.32 24.01 13.37 ;
      RECT 23.73 11.56 23.89 12.48 ;
      RECT 23.37 11.56 24.49 11.72 ;
      RECT 24.33 10.4 24.49 11.72 ;
      RECT 23.37 10.27 23.53 11.72 ;
      RECT 24.33 12 24.49 12.84 ;
      RECT 24.05 12 24.49 12.16 ;
      RECT 24.05 11.88 24.21 12.16 ;
      RECT 22.97 28.04 23.29 28.32 ;
      RECT 23.13 25.99 23.29 28.32 ;
      RECT 24.32 27.02 24.48 27.7 ;
      RECT 23.13 27.02 24.48 27.18 ;
      RECT 23.13 25.99 23.51 26.23 ;
      RECT 23.35 25.16 23.51 26.23 ;
      RECT 23.93 55.68 24.09 56.51 ;
      RECT 23.69 55.68 24.09 55.84 ;
      RECT 23.69 53.67 23.85 55.84 ;
      RECT 23.69 53.67 24.33 53.83 ;
      RECT 24.05 53.35 24.33 53.83 ;
      RECT 23.79 51.7 24.17 51.92 ;
      RECT 24.01 50.98 24.17 51.92 ;
      RECT 23.37 52.58 24.13 52.86 ;
      RECT 23.97 52.18 24.13 52.86 ;
      RECT 23.37 51.64 23.53 52.86 ;
      RECT 22.19 8.5 22.35 11.72 ;
      RECT 21.23 8.12 21.39 11.72 ;
      RECT 20.27 9.28 20.43 11.72 ;
      RECT 23.85 9.63 24.01 11.4 ;
      RECT 22.19 9.95 24.01 10.11 ;
      RECT 23.16 9.79 23.32 10.11 ;
      RECT 20.19 8.12 20.39 9.84 ;
      RECT 23.56 9.63 24.07 9.79 ;
      RECT 20.19 9.28 21.39 9.44 ;
      RECT 22.08 8.5 22.39 8.78 ;
      RECT 21.23 8.56 22.39 8.72 ;
      RECT 23.69 62.9 23.85 67.89 ;
      RECT 23.69 65.82 23.91 66.55 ;
      RECT 22.68 8.96 22.84 9.79 ;
      RECT 22.68 8.96 23.87 9.12 ;
      RECT 23.37 47.39 23.53 49.72 ;
      RECT 23.37 47.39 23.85 47.55 ;
      RECT 23.69 43.85 23.85 47.55 ;
      RECT 23.07 43.85 23.85 44.01 ;
      RECT 23.07 39.56 23.23 44.01 ;
      RECT 23.07 39.56 23.41 39.84 ;
      RECT 23.25 39.16 23.41 39.84 ;
      RECT 23.67 22.01 23.83 23.37 ;
      RECT 23.05 22.01 23.83 22.17 ;
      RECT 23.35 24.72 23.73 24.96 ;
      RECT 23.35 22.35 23.51 24.96 ;
      RECT 23.39 34.44 23.73 34.72 ;
      RECT 23.57 32.44 23.73 34.72 ;
      RECT 23.39 33.11 23.73 33.39 ;
      RECT 23.39 32.44 23.73 32.72 ;
      RECT 23.39 40.7 23.73 40.98 ;
      RECT 23.57 38.7 23.73 40.98 ;
      RECT 23.39 40.03 23.73 40.31 ;
      RECT 23.39 38.7 23.73 38.98 ;
      RECT 23.55 14.44 23.71 15.64 ;
      RECT 23.21 14.44 23.71 14.6 ;
      RECT 23.37 12.21 23.53 13.28 ;
      RECT 21.95 12.21 23.53 12.37 ;
      RECT 22.91 11.47 23.07 12.37 ;
      RECT 22.85 10.85 23.01 11.63 ;
      RECT 23.21 62.9 23.37 67.89 ;
      RECT 23.21 64.59 23.49 65.31 ;
      RECT 22.73 46.75 22.89 47.43 ;
      RECT 22.41 46.75 23.21 46.91 ;
      RECT 23.05 44.23 23.21 46.91 ;
      RECT 22.41 44.23 22.57 46.91 ;
      RECT 22.53 10.51 22.69 11.24 ;
      RECT 22.53 10.51 23.19 10.67 ;
      RECT 22.89 20.63 23.17 20.79 ;
      RECT 22.89 19.59 23.05 20.79 ;
      RECT 21.79 12.53 21.95 13.61 ;
      RECT 21.63 11.88 21.79 12.69 ;
      RECT 22.51 11.77 22.75 12.05 ;
      RECT 21.63 11.88 22.75 12.04 ;
      RECT 21.71 8.88 21.87 12.04 ;
      RECT 20.51 34.88 22.71 35.04 ;
      RECT 22.43 34.59 22.71 35.04 ;
      RECT 21.49 34.59 21.73 35.04 ;
      RECT 20.51 34.59 20.79 35.04 ;
      RECT 21.49 38.38 21.73 39.02 ;
      RECT 22.43 38.38 22.71 38.83 ;
      RECT 20.51 38.38 20.79 38.83 ;
      RECT 20.51 38.38 22.71 38.54 ;
      RECT 22.33 28.04 22.65 28.32 ;
      RECT 22.33 25.99 22.49 28.32 ;
      RECT 21.14 27.02 21.3 27.7 ;
      RECT 21.14 27.02 22.49 27.18 ;
      RECT 22.11 25.99 22.49 26.23 ;
      RECT 22.11 25.16 22.27 26.23 ;
      RECT 20.67 36.47 22.55 36.63 ;
      RECT 22.39 35.88 22.55 36.63 ;
      RECT 21.53 35.23 21.69 36.63 ;
      RECT 20.67 35.88 20.83 36.63 ;
      RECT 22.49 35.23 22.65 36.06 ;
      RECT 20.57 35.23 20.73 36.06 ;
      RECT 22.49 37.11 22.65 38.19 ;
      RECT 21.53 36.79 21.69 38.19 ;
      RECT 20.57 37.11 20.73 38.19 ;
      RECT 22.39 36.79 22.55 37.39 ;
      RECT 20.67 36.79 20.83 37.39 ;
      RECT 20.67 36.79 22.55 36.95 ;
      RECT 22.47 20.26 22.63 21.05 ;
      RECT 21.9 20.26 22.63 20.44 ;
      RECT 21.9 19.89 22.06 20.44 ;
      RECT 21.24 19.89 22.06 20.05 ;
      RECT 21.24 19.61 21.43 20.05 ;
      RECT 21.15 19.61 21.43 19.77 ;
      RECT 21.79 22.01 21.95 23.37 ;
      RECT 21.79 22.01 22.57 22.17 ;
      RECT 20.75 68.07 22.57 68.23 ;
      RECT 20.75 62.02 20.91 68.23 ;
      RECT 20.75 62.02 21.13 62.18 ;
      RECT 20.97 57.45 21.13 62.18 ;
      RECT 20.97 57.45 22.57 57.61 ;
      RECT 22.25 57.39 22.57 57.61 ;
      RECT 22.25 53.74 22.41 57.61 ;
      RECT 22.41 51.32 22.57 53.9 ;
      RECT 22.09 51.32 22.57 51.48 ;
      RECT 22.09 49.88 22.25 51.48 ;
      RECT 21.77 49.88 22.25 50.04 ;
      RECT 21.77 47.71 21.93 50.04 ;
      RECT 21.31 47.71 21.93 47.99 ;
      RECT 22.09 47.39 22.25 49.72 ;
      RECT 21.77 47.39 22.25 47.55 ;
      RECT 21.77 43.85 21.93 47.55 ;
      RECT 21.77 43.85 22.55 44.01 ;
      RECT 22.39 39.56 22.55 44.01 ;
      RECT 22.21 39.56 22.55 39.84 ;
      RECT 22.21 39.16 22.37 39.84 ;
      RECT 22.25 62.9 22.41 67.89 ;
      RECT 22.13 64.59 22.41 65.31 ;
      RECT 21.89 24.72 22.27 24.96 ;
      RECT 22.11 22.35 22.27 24.96 ;
      RECT 21.49 52.58 22.25 52.86 ;
      RECT 22.09 51.64 22.25 52.86 ;
      RECT 21.49 52.18 21.65 52.86 ;
      RECT 21.89 34.44 22.23 34.72 ;
      RECT 21.89 32.44 22.05 34.72 ;
      RECT 21.89 33.11 22.23 33.39 ;
      RECT 21.89 32.44 22.23 32.72 ;
      RECT 21.89 40.7 22.23 40.98 ;
      RECT 21.89 38.7 22.05 40.98 ;
      RECT 21.89 40.03 22.23 40.31 ;
      RECT 21.89 38.7 22.23 38.98 ;
      RECT 21.95 53.23 22.23 53.51 ;
      RECT 21.95 53.03 22.11 53.51 ;
      RECT 21.13 53.03 22.11 53.19 ;
      RECT 21.13 50.98 21.29 53.19 ;
      RECT 21.09 52.54 21.29 52.82 ;
      RECT 20.75 50.98 21.29 51.14 ;
      RECT 20.75 50.8 20.97 51.14 ;
      RECT 20.65 56.67 20.81 61.86 ;
      RECT 20.65 56.67 22.09 56.83 ;
      RECT 21.93 56 22.09 56.83 ;
      RECT 20.81 54.4 20.97 56.83 ;
      RECT 21.79 26.36 21.95 26.72 ;
      RECT 19.65 26.36 21.95 26.52 ;
      RECT 19.65 26.04 19.81 26.52 ;
      RECT 19 26.04 19.81 26.2 ;
      RECT 21.77 50.66 21.93 51.5 ;
      RECT 21.13 50.66 21.93 50.82 ;
      RECT 21.13 50.18 21.29 50.82 ;
      RECT 20.65 50.18 21.29 50.5 ;
      RECT 20.65 47.07 20.81 50.5 ;
      RECT 20.65 47.07 21.13 47.23 ;
      RECT 20.97 45.44 21.13 47.23 ;
      RECT 21.53 55.68 21.69 56.51 ;
      RECT 21.53 55.68 21.93 55.84 ;
      RECT 21.77 53.67 21.93 55.84 ;
      RECT 21.29 53.67 21.93 53.83 ;
      RECT 21.29 53.35 21.57 53.83 ;
      RECT 21.77 62.9 21.93 67.89 ;
      RECT 21.71 65.82 21.93 66.55 ;
      RECT 21.45 51.7 21.83 51.92 ;
      RECT 21.45 50.98 21.61 51.92 ;
      RECT 19.62 28.01 21.78 28.17 ;
      RECT 21.62 27.34 21.78 28.17 ;
      RECT 21.46 27.93 21.78 28.17 ;
      RECT 20.62 26.97 20.78 28.17 ;
      RECT 19.62 26.68 19.78 28.17 ;
      RECT 20.97 47.39 21.13 49.72 ;
      RECT 20.97 47.39 21.45 47.55 ;
      RECT 21.29 43.85 21.45 47.55 ;
      RECT 20.67 43.85 21.45 44.01 ;
      RECT 20.67 39.56 20.83 44.01 ;
      RECT 20.67 39.56 21.01 39.84 ;
      RECT 20.85 39.16 21.01 39.84 ;
      RECT 21.13 24.79 21.33 25.35 ;
      RECT 21.01 24.79 21.33 25.03 ;
      RECT 20.99 34.44 21.33 34.72 ;
      RECT 21.17 32.44 21.33 34.72 ;
      RECT 20.99 33.11 21.33 33.39 ;
      RECT 20.99 32.44 21.33 32.72 ;
      RECT 20.99 40.7 21.33 40.98 ;
      RECT 21.17 38.7 21.33 40.98 ;
      RECT 20.99 40.03 21.33 40.31 ;
      RECT 20.99 38.7 21.33 38.98 ;
      RECT 21.01 21.85 21.17 24.3 ;
      RECT 21.01 21.85 21.31 22.13 ;
      RECT 21.13 54.06 21.29 56.51 ;
      RECT 20.77 54.06 21.29 54.22 ;
      RECT 20.77 52.98 20.97 54.22 ;
      RECT 20.77 51.34 20.93 54.22 ;
      RECT 20.77 51.34 20.97 52.12 ;
      RECT 20.83 12.56 20.99 13.61 ;
      RECT 20.93 11.9 21.09 13.24 ;
      RECT 19.81 11.9 21.09 12.06 ;
      RECT 20.75 9.6 20.91 12.06 ;
      RECT 19.4 18.3 20.34 18.46 ;
      RECT 19.4 17.05 19.76 18.46 ;
      RECT 19.6 16.2 19.76 18.46 ;
      RECT 19.55 16.2 20.51 16.36 ;
      RECT 20.28 16.07 20.95 16.23 ;
      RECT 19.55 16.08 19.71 16.36 ;
      RECT 20.59 8.96 20.91 9.12 ;
      RECT 20.75 7.8 20.91 9.12 ;
      RECT 18.41 7.91 18.57 8.8 ;
      RECT 18.41 7.91 19.49 8.07 ;
      RECT 19.33 7.8 20.91 7.96 ;
      RECT 19.92 16.52 20.1 16.84 ;
      RECT 19.92 16.52 20.82 16.68 ;
      RECT 20.33 46.75 20.49 47.43 ;
      RECT 20.01 46.75 20.81 46.91 ;
      RECT 20.65 44.23 20.81 46.91 ;
      RECT 20.01 44.23 20.17 46.91 ;
      RECT 20.4 16.92 20.56 18.12 ;
      RECT 20.4 16.92 20.8 17.08 ;
      RECT 19.25 11.5 19.41 13.22 ;
      RECT 19.25 12.22 20.77 12.38 ;
      RECT 19.25 11.5 19.67 11.66 ;
      RECT 20.17 26.02 20.73 26.18 ;
      RECT 20.17 25.58 20.33 26.18 ;
      RECT 19.63 25.58 20.33 25.74 ;
      RECT 19.63 24 19.83 25.74 ;
      RECT 18.83 24.3 19.83 24.46 ;
      RECT 19.63 22.71 19.79 25.74 ;
      RECT 19.73 22.04 19.89 22.99 ;
      RECT 19.89 21.85 20.05 22.32 ;
      RECT 19.21 22.13 19.57 22.41 ;
      RECT 19.41 21.53 19.57 22.41 ;
      RECT 20.28 21.53 20.44 21.92 ;
      RECT 19.41 21.53 20.44 21.69 ;
      RECT 20.1 20.21 20.26 21.69 ;
      RECT 20.14 26.69 20.3 27.85 ;
      RECT 20.1 26.69 20.34 27.33 ;
      RECT 18.11 34.88 20.31 35.04 ;
      RECT 20.03 34.59 20.31 35.04 ;
      RECT 19.09 34.59 19.33 35.04 ;
      RECT 18.11 34.59 18.39 35.04 ;
      RECT 19.09 38.38 19.33 39.02 ;
      RECT 20.03 38.38 20.31 38.83 ;
      RECT 18.11 38.38 18.39 38.83 ;
      RECT 18.11 38.38 20.31 38.54 ;
      RECT 19.95 23.18 20.11 23.84 ;
      RECT 19.95 23.18 20.28 23.34 ;
      RECT 20.12 22.65 20.28 23.34 ;
      RECT 18.27 36.47 20.15 36.63 ;
      RECT 19.99 35.86 20.15 36.63 ;
      RECT 19.13 35.23 19.29 36.63 ;
      RECT 18.27 35.86 18.43 36.63 ;
      RECT 20.09 35.23 20.25 36.05 ;
      RECT 18.17 35.23 18.33 36.05 ;
      RECT 20.09 37.11 20.25 38.19 ;
      RECT 19.13 36.79 19.29 38.19 ;
      RECT 18.17 37.11 18.33 38.19 ;
      RECT 19.99 36.79 20.15 37.39 ;
      RECT 18.27 36.79 18.43 37.39 ;
      RECT 18.27 36.79 20.15 36.95 ;
      RECT 18.89 50.66 19.05 51.5 ;
      RECT 18.89 50.66 19.69 50.82 ;
      RECT 19.53 50.18 19.69 50.82 ;
      RECT 19.53 50.18 20.17 50.5 ;
      RECT 20.01 47.07 20.17 50.5 ;
      RECT 19.69 47.07 20.17 47.23 ;
      RECT 19.69 45.44 19.85 47.23 ;
      RECT 20.01 56.67 20.17 61.86 ;
      RECT 18.73 56.67 20.17 56.83 ;
      RECT 19.85 54.4 20.01 56.83 ;
      RECT 18.73 56 18.89 56.83 ;
      RECT 19.69 47.39 19.85 49.72 ;
      RECT 19.37 47.39 19.85 47.55 ;
      RECT 19.37 43.85 19.53 47.55 ;
      RECT 19.37 43.85 20.15 44.01 ;
      RECT 19.99 39.56 20.15 44.01 ;
      RECT 19.81 39.56 20.15 39.84 ;
      RECT 19.81 39.16 19.97 39.84 ;
      RECT 18.6 28.52 19.69 28.68 ;
      RECT 19.41 28.35 19.69 28.68 ;
      RECT 19.41 28.35 20.09 28.51 ;
      RECT 18.59 53.23 18.87 53.51 ;
      RECT 18.71 53.03 18.87 53.51 ;
      RECT 18.71 53.03 19.69 53.19 ;
      RECT 19.53 50.98 19.69 53.19 ;
      RECT 19.53 52.54 19.73 52.82 ;
      RECT 19.53 50.98 20.07 51.14 ;
      RECT 19.85 50.8 20.07 51.14 ;
      RECT 18.25 68.07 20.07 68.23 ;
      RECT 19.91 62.02 20.07 68.23 ;
      RECT 19.69 62.02 20.07 62.18 ;
      RECT 19.69 57.45 19.85 62.18 ;
      RECT 18.25 57.45 19.85 57.61 ;
      RECT 18.25 57.39 18.57 57.61 ;
      RECT 18.41 53.74 18.57 57.61 ;
      RECT 18.25 51.32 18.41 53.9 ;
      RECT 18.25 51.32 18.73 51.48 ;
      RECT 18.57 49.88 18.73 51.48 ;
      RECT 18.57 49.88 19.05 50.04 ;
      RECT 18.89 47.71 19.05 50.04 ;
      RECT 18.89 47.71 19.51 47.99 ;
      RECT 19.53 54.06 19.69 56.51 ;
      RECT 19.53 54.06 20.05 54.22 ;
      RECT 19.89 51.34 20.05 54.22 ;
      RECT 19.85 52.98 20.05 54.22 ;
      RECT 19.85 51.34 20.05 52.12 ;
      RECT 18.73 12.92 18.89 13.67 ;
      RECT 18.73 12.92 19.09 13.08 ;
      RECT 18.93 9.68 19.09 13.08 ;
      RECT 18.89 9.68 19.09 11.89 ;
      RECT 18.89 9.68 19.87 9.84 ;
      RECT 19.71 8.6 19.87 9.84 ;
      RECT 19.49 34.44 19.83 34.72 ;
      RECT 19.49 32.44 19.65 34.72 ;
      RECT 19.49 33.11 19.83 33.39 ;
      RECT 19.49 32.44 19.83 32.72 ;
      RECT 19.49 40.7 19.83 40.98 ;
      RECT 19.49 38.7 19.65 40.98 ;
      RECT 19.49 40.03 19.83 40.31 ;
      RECT 19.49 38.7 19.83 38.98 ;
      RECT 19.13 55.68 19.29 56.51 ;
      RECT 18.89 55.68 19.29 55.84 ;
      RECT 18.89 53.67 19.05 55.84 ;
      RECT 18.89 53.67 19.53 53.83 ;
      RECT 19.25 53.35 19.53 53.83 ;
      RECT 19.08 16.52 19.24 18.9 ;
      RECT 19.08 16.52 19.44 16.8 ;
      RECT 19.21 15.31 19.37 16.8 ;
      RECT 18.68 24.79 18.84 28.32 ;
      RECT 18.68 25.16 19.37 25.32 ;
      RECT 18.99 51.7 19.37 51.92 ;
      RECT 19.21 50.98 19.37 51.92 ;
      RECT 18.57 52.58 19.33 52.86 ;
      RECT 19.17 52.18 19.33 52.86 ;
      RECT 18.57 51.64 18.73 52.86 ;
      RECT 18.41 23.98 18.59 24.52 ;
      RECT 18.41 23.98 19.11 24.14 ;
      RECT 18.95 23.27 19.11 24.14 ;
      RECT 18.89 21.78 19.05 23.43 ;
      RECT 19.03 21.21 19.19 21.94 ;
      RECT 19.16 20.95 19.32 21.37 ;
      RECT 17.93 7.5 18.09 8.72 ;
      RECT 17.93 7.58 18.14 7.9 ;
      RECT 17.93 7.59 19.17 7.75 ;
      RECT 17.93 7.58 18.21 7.75 ;
      RECT 18.89 62.9 19.05 67.89 ;
      RECT 18.89 65.82 19.11 66.55 ;
      RECT 18.57 47.39 18.73 49.72 ;
      RECT 18.57 47.39 19.05 47.55 ;
      RECT 18.89 43.85 19.05 47.55 ;
      RECT 18.27 43.85 19.05 44.01 ;
      RECT 18.27 39.56 18.43 44.01 ;
      RECT 18.27 39.56 18.61 39.84 ;
      RECT 18.45 39.16 18.61 39.84 ;
      RECT 18.59 34.44 18.93 34.72 ;
      RECT 18.77 32.44 18.93 34.72 ;
      RECT 18.59 33.11 18.93 33.39 ;
      RECT 18.59 32.44 18.93 32.72 ;
      RECT 18.59 40.7 18.93 40.98 ;
      RECT 18.77 38.7 18.93 40.98 ;
      RECT 18.59 40.03 18.93 40.31 ;
      RECT 18.59 38.7 18.93 38.98 ;
      RECT 18.16 15.57 18.32 17.28 ;
      RECT 18.76 16.43 18.92 16.71 ;
      RECT 18.16 16.43 18.92 16.59 ;
      RECT 18.1 15.57 18.38 15.73 ;
      RECT 18.6 17.18 18.76 18.9 ;
      RECT 17.93 17.96 18.76 18.12 ;
      RECT 17.93 17.84 18.09 18.12 ;
      RECT 18.64 17.06 18.8 17.34 ;
      RECT 18.25 23.66 18.79 23.82 ;
      RECT 18.25 20.12 18.41 23.82 ;
      RECT 18.25 23.22 18.71 23.38 ;
      RECT 18.16 20.83 18.41 21.11 ;
      RECT 18.25 20.12 18.68 20.28 ;
      RECT 18.41 62.9 18.57 67.89 ;
      RECT 18.41 64.59 18.69 65.31 ;
      RECT 18.45 10.08 18.61 11.89 ;
      RECT 17.87 10.08 18.61 10.24 ;
      RECT 17.93 8.88 18.09 10.24 ;
      RECT 17.93 46.75 18.09 47.43 ;
      RECT 17.61 46.75 18.41 46.91 ;
      RECT 18.25 44.23 18.41 46.91 ;
      RECT 17.61 44.23 17.77 46.91 ;
      RECT 18.2 26.15 18.36 28.96 ;
      RECT 18.17 26.15 18.36 26.51 ;
      RECT 15.71 34.88 17.91 35.04 ;
      RECT 17.63 34.59 17.91 35.04 ;
      RECT 16.69 34.59 16.93 35.04 ;
      RECT 15.71 34.59 15.99 35.04 ;
      RECT 16.69 38.38 16.93 39.02 ;
      RECT 17.63 38.38 17.91 38.83 ;
      RECT 15.71 38.38 15.99 38.83 ;
      RECT 15.71 38.38 17.91 38.54 ;
      RECT 15.87 36.47 17.75 36.63 ;
      RECT 17.59 35.88 17.75 36.63 ;
      RECT 16.73 35.23 16.89 36.63 ;
      RECT 15.87 35.88 16.03 36.63 ;
      RECT 17.69 35.23 17.85 36.06 ;
      RECT 15.77 35.23 15.93 36.06 ;
      RECT 17.69 37.11 17.85 38.19 ;
      RECT 16.73 36.79 16.89 38.19 ;
      RECT 15.77 37.11 15.93 38.19 ;
      RECT 17.59 36.79 17.75 37.39 ;
      RECT 15.87 36.79 16.03 37.39 ;
      RECT 15.87 36.79 17.75 36.95 ;
      RECT 15.95 68.07 17.77 68.23 ;
      RECT 15.95 62.02 16.11 68.23 ;
      RECT 15.95 62.02 16.33 62.18 ;
      RECT 16.17 57.45 16.33 62.18 ;
      RECT 16.17 57.45 17.77 57.61 ;
      RECT 17.45 57.39 17.77 57.61 ;
      RECT 17.45 53.74 17.61 57.61 ;
      RECT 17.61 51.32 17.77 53.9 ;
      RECT 17.29 51.32 17.77 51.48 ;
      RECT 17.29 49.88 17.45 51.48 ;
      RECT 16.97 49.88 17.45 50.04 ;
      RECT 16.97 47.71 17.13 50.04 ;
      RECT 16.51 47.71 17.13 47.99 ;
      RECT 17.29 47.39 17.45 49.72 ;
      RECT 16.97 47.39 17.45 47.55 ;
      RECT 16.97 43.85 17.13 47.55 ;
      RECT 16.97 43.85 17.75 44.01 ;
      RECT 17.59 39.56 17.75 44.01 ;
      RECT 17.41 39.56 17.75 39.84 ;
      RECT 17.41 39.16 17.57 39.84 ;
      RECT 17.45 62.9 17.61 67.89 ;
      RECT 17.33 64.59 17.61 65.31 ;
      RECT 16.69 52.58 17.45 52.86 ;
      RECT 17.29 51.64 17.45 52.86 ;
      RECT 16.69 52.18 16.85 52.86 ;
      RECT 17.09 34.44 17.43 34.72 ;
      RECT 17.09 32.44 17.25 34.72 ;
      RECT 17.09 33.11 17.43 33.39 ;
      RECT 17.09 32.44 17.43 32.72 ;
      RECT 17.09 40.7 17.43 40.98 ;
      RECT 17.09 38.7 17.25 40.98 ;
      RECT 17.09 40.03 17.43 40.31 ;
      RECT 17.09 38.7 17.43 38.98 ;
      RECT 17.15 53.23 17.43 53.51 ;
      RECT 17.15 53.03 17.31 53.51 ;
      RECT 16.33 53.03 17.31 53.19 ;
      RECT 16.33 50.98 16.49 53.19 ;
      RECT 16.29 52.54 16.49 52.82 ;
      RECT 15.95 50.98 16.49 51.14 ;
      RECT 15.95 50.8 16.17 51.14 ;
      RECT 15.85 56.67 16.01 61.86 ;
      RECT 15.85 56.67 17.29 56.83 ;
      RECT 17.13 56 17.29 56.83 ;
      RECT 16.01 54.4 16.17 56.83 ;
      RECT 9.29 12.95 17.13 13.55 ;
      RECT 16.53 8.34 17.13 13.55 ;
      RECT 9.29 8.34 9.89 13.55 ;
      RECT 9.29 8.34 17.13 8.88 ;
      RECT 9.29 26.87 17.13 27.47 ;
      RECT 16.53 18.71 17.13 27.47 ;
      RECT 9.29 18.71 9.89 27.47 ;
      RECT 9.29 24.41 17.13 25.01 ;
      RECT 9.29 18.71 17.13 19.31 ;
      RECT 16.97 50.66 17.13 51.5 ;
      RECT 16.33 50.66 17.13 50.82 ;
      RECT 16.33 50.18 16.49 50.82 ;
      RECT 15.85 50.18 16.49 50.5 ;
      RECT 15.85 47.07 16.01 50.5 ;
      RECT 15.85 47.07 16.33 47.23 ;
      RECT 16.17 45.44 16.33 47.23 ;
      RECT 16.73 55.68 16.89 56.51 ;
      RECT 16.73 55.68 17.13 55.84 ;
      RECT 16.97 53.67 17.13 55.84 ;
      RECT 16.49 53.67 17.13 53.83 ;
      RECT 16.49 53.35 16.77 53.83 ;
      RECT 16.97 62.9 17.13 67.89 ;
      RECT 16.91 65.82 17.13 66.55 ;
      RECT 16.65 51.7 17.03 51.92 ;
      RECT 16.65 50.98 16.81 51.92 ;
      RECT 16.17 47.39 16.33 49.72 ;
      RECT 16.17 47.39 16.65 47.55 ;
      RECT 16.49 43.85 16.65 47.55 ;
      RECT 15.87 43.85 16.65 44.01 ;
      RECT 15.87 39.56 16.03 44.01 ;
      RECT 15.87 39.56 16.21 39.84 ;
      RECT 16.05 39.16 16.21 39.84 ;
      RECT 16.19 34.44 16.53 34.72 ;
      RECT 16.37 32.44 16.53 34.72 ;
      RECT 16.19 33.11 16.53 33.39 ;
      RECT 16.19 32.44 16.53 32.72 ;
      RECT 16.19 40.7 16.53 40.98 ;
      RECT 16.37 38.7 16.53 40.98 ;
      RECT 16.19 40.03 16.53 40.31 ;
      RECT 16.19 38.7 16.53 38.98 ;
      RECT 16.33 54.06 16.49 56.51 ;
      RECT 15.97 54.06 16.49 54.22 ;
      RECT 15.97 52.98 16.17 54.22 ;
      RECT 15.97 51.34 16.13 54.22 ;
      RECT 15.97 51.34 16.17 52.12 ;
      RECT 15.53 46.75 15.69 47.43 ;
      RECT 15.21 46.75 16.01 46.91 ;
      RECT 15.85 44.23 16.01 46.91 ;
      RECT 15.21 44.23 15.37 46.91 ;
      RECT 13.31 34.88 15.51 35.04 ;
      RECT 15.23 34.59 15.51 35.04 ;
      RECT 14.29 34.59 14.53 35.04 ;
      RECT 13.31 34.59 13.59 35.04 ;
      RECT 14.29 38.38 14.53 39.02 ;
      RECT 15.23 38.38 15.51 38.83 ;
      RECT 13.31 38.38 13.59 38.83 ;
      RECT 13.31 38.38 15.51 38.54 ;
      RECT 13.47 36.47 15.35 36.63 ;
      RECT 15.19 35.86 15.35 36.63 ;
      RECT 14.33 35.23 14.49 36.63 ;
      RECT 13.47 35.86 13.63 36.63 ;
      RECT 15.29 35.23 15.45 36.05 ;
      RECT 13.37 35.23 13.53 36.05 ;
      RECT 15.29 37.11 15.45 38.19 ;
      RECT 14.33 36.79 14.49 38.19 ;
      RECT 13.37 37.11 13.53 38.19 ;
      RECT 15.19 36.79 15.35 37.39 ;
      RECT 13.47 36.79 13.63 37.39 ;
      RECT 13.47 36.79 15.35 36.95 ;
      RECT 14.09 50.66 14.25 51.5 ;
      RECT 14.09 50.66 14.89 50.82 ;
      RECT 14.73 50.18 14.89 50.82 ;
      RECT 14.73 50.18 15.37 50.5 ;
      RECT 15.21 47.07 15.37 50.5 ;
      RECT 14.89 47.07 15.37 47.23 ;
      RECT 14.89 45.44 15.05 47.23 ;
      RECT 15.21 56.67 15.37 61.86 ;
      RECT 13.93 56.67 15.37 56.83 ;
      RECT 15.05 54.4 15.21 56.83 ;
      RECT 13.93 56 14.09 56.83 ;
      RECT 14.89 47.39 15.05 49.72 ;
      RECT 14.57 47.39 15.05 47.55 ;
      RECT 14.57 43.85 14.73 47.55 ;
      RECT 14.57 43.85 15.35 44.01 ;
      RECT 15.19 39.56 15.35 44.01 ;
      RECT 15.01 39.56 15.35 39.84 ;
      RECT 15.01 39.16 15.17 39.84 ;
      RECT 13.79 53.23 14.07 53.51 ;
      RECT 13.91 53.03 14.07 53.51 ;
      RECT 13.91 53.03 14.89 53.19 ;
      RECT 14.73 50.98 14.89 53.19 ;
      RECT 14.73 52.54 14.93 52.82 ;
      RECT 14.73 50.98 15.27 51.14 ;
      RECT 15.05 50.8 15.27 51.14 ;
      RECT 13.45 68.07 15.27 68.23 ;
      RECT 15.11 62.02 15.27 68.23 ;
      RECT 14.89 62.02 15.27 62.18 ;
      RECT 14.89 57.45 15.05 62.18 ;
      RECT 13.45 57.45 15.05 57.61 ;
      RECT 13.45 57.39 13.77 57.61 ;
      RECT 13.61 53.74 13.77 57.61 ;
      RECT 13.45 51.32 13.61 53.9 ;
      RECT 13.45 51.32 13.93 51.48 ;
      RECT 13.77 49.88 13.93 51.48 ;
      RECT 13.77 49.88 14.25 50.04 ;
      RECT 14.09 47.71 14.25 50.04 ;
      RECT 14.09 47.71 14.71 47.99 ;
      RECT 14.73 54.06 14.89 56.51 ;
      RECT 14.73 54.06 15.25 54.22 ;
      RECT 15.09 51.34 15.25 54.22 ;
      RECT 15.05 52.98 15.25 54.22 ;
      RECT 15.05 51.34 15.25 52.12 ;
      RECT 14.69 34.44 15.03 34.72 ;
      RECT 14.69 32.44 14.85 34.72 ;
      RECT 14.69 33.11 15.03 33.39 ;
      RECT 14.69 32.44 15.03 32.72 ;
      RECT 14.69 40.7 15.03 40.98 ;
      RECT 14.69 38.7 14.85 40.98 ;
      RECT 14.69 40.03 15.03 40.31 ;
      RECT 14.69 38.7 15.03 38.98 ;
      RECT 14.33 55.68 14.49 56.51 ;
      RECT 14.09 55.68 14.49 55.84 ;
      RECT 14.09 53.67 14.25 55.84 ;
      RECT 14.09 53.67 14.73 53.83 ;
      RECT 14.45 53.35 14.73 53.83 ;
      RECT 14.19 51.7 14.57 51.92 ;
      RECT 14.41 50.98 14.57 51.92 ;
      RECT 13.77 52.58 14.53 52.86 ;
      RECT 14.37 52.18 14.53 52.86 ;
      RECT 13.77 51.64 13.93 52.86 ;
      RECT 14.09 62.9 14.25 67.89 ;
      RECT 14.09 65.82 14.31 66.55 ;
      RECT 13.77 47.39 13.93 49.72 ;
      RECT 13.77 47.39 14.25 47.55 ;
      RECT 14.09 43.85 14.25 47.55 ;
      RECT 13.47 43.85 14.25 44.01 ;
      RECT 13.47 39.56 13.63 44.01 ;
      RECT 13.47 39.56 13.81 39.84 ;
      RECT 13.65 39.16 13.81 39.84 ;
      RECT 13.79 34.44 14.13 34.72 ;
      RECT 13.97 32.44 14.13 34.72 ;
      RECT 13.79 33.11 14.13 33.39 ;
      RECT 13.79 32.44 14.13 32.72 ;
      RECT 13.79 40.7 14.13 40.98 ;
      RECT 13.97 38.7 14.13 40.98 ;
      RECT 13.79 40.03 14.13 40.31 ;
      RECT 13.79 38.7 14.13 38.98 ;
      RECT 13.61 62.9 13.77 67.89 ;
      RECT 13.61 64.59 13.89 65.31 ;
      RECT 13.13 46.75 13.29 47.43 ;
      RECT 12.81 46.75 13.61 46.91 ;
      RECT 13.45 44.23 13.61 46.91 ;
      RECT 12.81 44.23 12.97 46.91 ;
      RECT 10.91 34.88 13.11 35.04 ;
      RECT 12.83 34.59 13.11 35.04 ;
      RECT 11.89 34.59 12.13 35.04 ;
      RECT 10.91 34.59 11.19 35.04 ;
      RECT 11.89 38.38 12.13 39.02 ;
      RECT 12.83 38.38 13.11 38.83 ;
      RECT 10.91 38.38 11.19 38.83 ;
      RECT 10.91 38.38 13.11 38.54 ;
      RECT 11.07 36.47 12.95 36.63 ;
      RECT 12.79 35.88 12.95 36.63 ;
      RECT 11.93 35.23 12.09 36.63 ;
      RECT 11.07 35.88 11.23 36.63 ;
      RECT 12.89 35.23 13.05 36.06 ;
      RECT 10.97 35.23 11.13 36.06 ;
      RECT 12.89 37.11 13.05 38.19 ;
      RECT 11.93 36.79 12.09 38.19 ;
      RECT 10.97 37.11 11.13 38.19 ;
      RECT 12.79 36.79 12.95 37.39 ;
      RECT 11.07 36.79 11.23 37.39 ;
      RECT 11.07 36.79 12.95 36.95 ;
      RECT 11.15 68.07 12.97 68.23 ;
      RECT 11.15 62.02 11.31 68.23 ;
      RECT 11.15 62.02 11.53 62.18 ;
      RECT 11.37 57.45 11.53 62.18 ;
      RECT 11.37 57.45 12.97 57.61 ;
      RECT 12.65 57.39 12.97 57.61 ;
      RECT 12.65 53.74 12.81 57.61 ;
      RECT 12.81 51.32 12.97 53.9 ;
      RECT 12.49 51.32 12.97 51.48 ;
      RECT 12.49 49.88 12.65 51.48 ;
      RECT 12.17 49.88 12.65 50.04 ;
      RECT 12.17 47.71 12.33 50.04 ;
      RECT 11.71 47.71 12.33 47.99 ;
      RECT 12.49 47.39 12.65 49.72 ;
      RECT 12.17 47.39 12.65 47.55 ;
      RECT 12.17 43.85 12.33 47.55 ;
      RECT 12.17 43.85 12.95 44.01 ;
      RECT 12.79 39.56 12.95 44.01 ;
      RECT 12.61 39.56 12.95 39.84 ;
      RECT 12.61 39.16 12.77 39.84 ;
      RECT 12.65 62.9 12.81 67.89 ;
      RECT 12.53 64.59 12.81 65.31 ;
      RECT 11.89 52.58 12.65 52.86 ;
      RECT 12.49 51.64 12.65 52.86 ;
      RECT 11.89 52.18 12.05 52.86 ;
      RECT 12.29 34.44 12.63 34.72 ;
      RECT 12.29 32.44 12.45 34.72 ;
      RECT 12.29 33.11 12.63 33.39 ;
      RECT 12.29 32.44 12.63 32.72 ;
      RECT 12.29 40.7 12.63 40.98 ;
      RECT 12.29 38.7 12.45 40.98 ;
      RECT 12.29 40.03 12.63 40.31 ;
      RECT 12.29 38.7 12.63 38.98 ;
      RECT 12.35 53.23 12.63 53.51 ;
      RECT 12.35 53.03 12.51 53.51 ;
      RECT 11.53 53.03 12.51 53.19 ;
      RECT 11.53 50.98 11.69 53.19 ;
      RECT 11.49 52.54 11.69 52.82 ;
      RECT 11.15 50.98 11.69 51.14 ;
      RECT 11.15 50.8 11.37 51.14 ;
      RECT 11.05 56.67 11.21 61.86 ;
      RECT 11.05 56.67 12.49 56.83 ;
      RECT 12.33 56 12.49 56.83 ;
      RECT 11.21 54.4 11.37 56.83 ;
      RECT 12.17 50.66 12.33 51.5 ;
      RECT 11.53 50.66 12.33 50.82 ;
      RECT 11.53 50.18 11.69 50.82 ;
      RECT 11.05 50.18 11.69 50.5 ;
      RECT 11.05 47.07 11.21 50.5 ;
      RECT 11.05 47.07 11.53 47.23 ;
      RECT 11.37 45.44 11.53 47.23 ;
      RECT 11.93 55.68 12.09 56.51 ;
      RECT 11.93 55.68 12.33 55.84 ;
      RECT 12.17 53.67 12.33 55.84 ;
      RECT 11.69 53.67 12.33 53.83 ;
      RECT 11.69 53.35 11.97 53.83 ;
      RECT 12.17 62.9 12.33 67.89 ;
      RECT 12.11 65.82 12.33 66.55 ;
      RECT 11.85 51.7 12.23 51.92 ;
      RECT 11.85 50.98 12.01 51.92 ;
      RECT 11.37 47.39 11.53 49.72 ;
      RECT 11.37 47.39 11.85 47.55 ;
      RECT 11.69 43.85 11.85 47.55 ;
      RECT 11.07 43.85 11.85 44.01 ;
      RECT 11.07 39.56 11.23 44.01 ;
      RECT 11.07 39.56 11.41 39.84 ;
      RECT 11.25 39.16 11.41 39.84 ;
      RECT 11.39 34.44 11.73 34.72 ;
      RECT 11.57 32.44 11.73 34.72 ;
      RECT 11.39 33.11 11.73 33.39 ;
      RECT 11.39 32.44 11.73 32.72 ;
      RECT 11.39 40.7 11.73 40.98 ;
      RECT 11.57 38.7 11.73 40.98 ;
      RECT 11.39 40.03 11.73 40.31 ;
      RECT 11.39 38.7 11.73 38.98 ;
      RECT 11.53 54.06 11.69 56.51 ;
      RECT 11.17 54.06 11.69 54.22 ;
      RECT 11.17 52.98 11.37 54.22 ;
      RECT 11.17 51.34 11.33 54.22 ;
      RECT 11.17 51.34 11.37 52.12 ;
      RECT 10.73 46.75 10.89 47.43 ;
      RECT 10.41 46.75 11.21 46.91 ;
      RECT 11.05 44.23 11.21 46.91 ;
      RECT 10.41 44.23 10.57 46.91 ;
      RECT 8.51 34.88 10.71 35.04 ;
      RECT 10.43 34.59 10.71 35.04 ;
      RECT 9.49 34.59 9.73 35.04 ;
      RECT 8.51 34.59 8.79 35.04 ;
      RECT 9.49 38.38 9.73 39.02 ;
      RECT 10.43 38.38 10.71 38.83 ;
      RECT 8.51 38.38 8.79 38.83 ;
      RECT 8.51 38.38 10.71 38.54 ;
      RECT 8.67 36.47 10.55 36.63 ;
      RECT 10.39 35.86 10.55 36.63 ;
      RECT 9.53 35.23 9.69 36.63 ;
      RECT 8.67 35.86 8.83 36.63 ;
      RECT 10.49 35.23 10.65 36.05 ;
      RECT 8.57 35.23 8.73 36.05 ;
      RECT 10.49 37.11 10.65 38.19 ;
      RECT 9.53 36.79 9.69 38.19 ;
      RECT 8.57 37.11 8.73 38.19 ;
      RECT 10.39 36.79 10.55 37.39 ;
      RECT 8.67 36.79 8.83 37.39 ;
      RECT 8.67 36.79 10.55 36.95 ;
      RECT 9.29 50.66 9.45 51.5 ;
      RECT 9.29 50.66 10.09 50.82 ;
      RECT 9.93 50.18 10.09 50.82 ;
      RECT 9.93 50.18 10.57 50.5 ;
      RECT 10.41 47.07 10.57 50.5 ;
      RECT 10.09 47.07 10.57 47.23 ;
      RECT 10.09 45.44 10.25 47.23 ;
      RECT 10.41 56.67 10.57 61.86 ;
      RECT 9.13 56.67 10.57 56.83 ;
      RECT 10.25 54.4 10.41 56.83 ;
      RECT 9.13 56 9.29 56.83 ;
      RECT 10.09 47.39 10.25 49.72 ;
      RECT 9.77 47.39 10.25 47.55 ;
      RECT 9.77 43.85 9.93 47.55 ;
      RECT 9.77 43.85 10.55 44.01 ;
      RECT 10.39 39.56 10.55 44.01 ;
      RECT 10.21 39.56 10.55 39.84 ;
      RECT 10.21 39.16 10.37 39.84 ;
      RECT 8.99 53.23 9.27 53.51 ;
      RECT 9.11 53.03 9.27 53.51 ;
      RECT 9.11 53.03 10.09 53.19 ;
      RECT 9.93 50.98 10.09 53.19 ;
      RECT 9.93 52.54 10.13 52.82 ;
      RECT 9.93 50.98 10.47 51.14 ;
      RECT 10.25 50.8 10.47 51.14 ;
      RECT 8.65 68.07 10.47 68.23 ;
      RECT 10.31 62.02 10.47 68.23 ;
      RECT 10.09 62.02 10.47 62.18 ;
      RECT 10.09 57.45 10.25 62.18 ;
      RECT 8.65 57.45 10.25 57.61 ;
      RECT 8.65 57.39 8.97 57.61 ;
      RECT 8.81 53.74 8.97 57.61 ;
      RECT 8.65 51.32 8.81 53.9 ;
      RECT 8.65 51.32 9.13 51.48 ;
      RECT 8.97 49.88 9.13 51.48 ;
      RECT 8.97 49.88 9.45 50.04 ;
      RECT 9.29 47.71 9.45 50.04 ;
      RECT 9.29 47.71 9.91 47.99 ;
      RECT 9.93 54.06 10.09 56.51 ;
      RECT 9.93 54.06 10.45 54.22 ;
      RECT 10.29 51.34 10.45 54.22 ;
      RECT 10.25 52.98 10.45 54.22 ;
      RECT 10.25 51.34 10.45 52.12 ;
      RECT 9.89 34.44 10.23 34.72 ;
      RECT 9.89 32.44 10.05 34.72 ;
      RECT 9.89 33.11 10.23 33.39 ;
      RECT 9.89 32.44 10.23 32.72 ;
      RECT 9.89 40.7 10.23 40.98 ;
      RECT 9.89 38.7 10.05 40.98 ;
      RECT 9.89 40.03 10.23 40.31 ;
      RECT 9.89 38.7 10.23 38.98 ;
      RECT 9.53 55.68 9.69 56.51 ;
      RECT 9.29 55.68 9.69 55.84 ;
      RECT 9.29 53.67 9.45 55.84 ;
      RECT 9.29 53.67 9.93 53.83 ;
      RECT 9.65 53.35 9.93 53.83 ;
      RECT 9.39 51.7 9.77 51.92 ;
      RECT 9.61 50.98 9.77 51.92 ;
      RECT 8.97 52.58 9.73 52.86 ;
      RECT 9.57 52.18 9.73 52.86 ;
      RECT 8.97 51.64 9.13 52.86 ;
      RECT 9.29 62.9 9.45 67.89 ;
      RECT 9.29 65.82 9.51 66.55 ;
      RECT 8.97 47.39 9.13 49.72 ;
      RECT 8.97 47.39 9.45 47.55 ;
      RECT 9.29 43.85 9.45 47.55 ;
      RECT 8.67 43.85 9.45 44.01 ;
      RECT 8.67 39.56 8.83 44.01 ;
      RECT 8.67 39.56 9.01 39.84 ;
      RECT 8.85 39.16 9.01 39.84 ;
      RECT 8.99 34.44 9.33 34.72 ;
      RECT 9.17 32.44 9.33 34.72 ;
      RECT 8.99 33.11 9.33 33.39 ;
      RECT 8.99 32.44 9.33 32.72 ;
      RECT 8.99 40.7 9.33 40.98 ;
      RECT 9.17 38.7 9.33 40.98 ;
      RECT 8.99 40.03 9.33 40.31 ;
      RECT 8.99 38.7 9.33 38.98 ;
      RECT 8.81 62.9 8.97 67.89 ;
      RECT 8.81 64.59 9.09 65.31 ;
      RECT 8.33 46.75 8.49 47.43 ;
      RECT 8.33 46.75 8.81 46.91 ;
      RECT 8.65 44.23 8.81 46.91 ;
      RECT 233.78 7.94 234.36 9.14 ;
      RECT 233.78 17.26 234.36 18.46 ;
      RECT 233.78 25.81 234.36 27.81 ;
      RECT 233.78 35.91 234.36 36.91 ;
      RECT 233.78 50.24 234.36 51.24 ;
      RECT 233.78 57.02 234.36 58.02 ;
      RECT 233.78 60.6 234.36 61.6 ;
      RECT 233.78 62.45 234.36 63.45 ;
      RECT 233.78 69.16 234.36 69.96 ;
      RECT 233.78 72.56 234.36 73.36 ;
      RECT 233.78 75.96 234.36 76.76 ;
      RECT 233.78 79.36 234.36 80.16 ;
      RECT 233.78 82.76 234.36 83.56 ;
      RECT 233.78 86.16 234.36 86.96 ;
      RECT 233.78 89.56 234.36 90.36 ;
      RECT 233.78 92.96 234.36 93.76 ;
      RECT 233.78 96.36 234.36 97.16 ;
      RECT 233.78 99.76 234.36 100.56 ;
      RECT 233.78 103.16 234.36 103.96 ;
      RECT 233.78 106.56 234.36 107.36 ;
      RECT 233.78 109.96 234.36 110.76 ;
      RECT 233.78 113.36 234.36 114.16 ;
      RECT 233.78 116.76 234.36 117.56 ;
      RECT 233.78 120.16 234.36 120.96 ;
      RECT 233.78 123.56 234.36 124.36 ;
      RECT 233.78 126.96 234.36 127.76 ;
      RECT 233.78 130.36 234.36 131.16 ;
      RECT 233.78 133.76 234.36 134.56 ;
      RECT 233.78 137.16 234.36 137.96 ;
      RECT 233.78 140.56 234.36 141.36 ;
      RECT 233.78 143.96 234.36 144.76 ;
      RECT 233.78 147.36 234.36 148.16 ;
      RECT 233.78 150.76 234.36 151.56 ;
      RECT 233.78 154.16 234.36 154.96 ;
      RECT 233.78 157.56 234.36 158.36 ;
      RECT 233.78 160.96 234.36 161.76 ;
      RECT 233.78 164.36 234.36 165.16 ;
      RECT 233.78 167.76 234.36 168.56 ;
      RECT 233.78 171.16 234.36 171.96 ;
      RECT 233.78 174.56 234.36 175.36 ;
      RECT 233.78 177.96 234.36 178.76 ;
      RECT 233.78 181.36 234.36 182.16 ;
      RECT 233.78 184.76 234.36 185.56 ;
      RECT 233.78 188.16 234.36 188.96 ;
      RECT 233.78 191.56 234.36 192.36 ;
      RECT 233.78 194.96 234.36 195.76 ;
      RECT 233.78 198.36 234.36 199.16 ;
      RECT 233.78 201.76 234.36 202.56 ;
      RECT 233.78 205.16 234.36 205.96 ;
      RECT 233.78 208.56 234.36 209.36 ;
      RECT 233.78 211.96 234.36 212.76 ;
      RECT 233.78 215.36 234.36 216.16 ;
      RECT 233.78 218.76 234.36 219.56 ;
      RECT 233.78 222.16 234.36 222.96 ;
      RECT 233.78 225.56 234.36 226.36 ;
      RECT 233.78 228.96 234.36 229.76 ;
      RECT 233.78 232.36 234.36 233.16 ;
      RECT 233.78 235.76 234.36 236.56 ;
      RECT 233.78 239.16 234.36 239.96 ;
      RECT 233.78 242.56 234.36 243.36 ;
      RECT 233.78 245.96 234.36 246.76 ;
      RECT 233.78 249.36 234.36 250.16 ;
      RECT 233.78 252.76 234.36 253.56 ;
      RECT 233.78 256.16 234.36 256.96 ;
      RECT 233.78 259.56 234.36 260.36 ;
      RECT 233.78 262.96 234.36 263.76 ;
      RECT 233.78 266.36 234.36 267.16 ;
      RECT 233.78 269.76 234.36 270.56 ;
      RECT 233.78 273.16 234.36 273.96 ;
      RECT 233.78 276.56 234.36 277.36 ;
      RECT 233.78 279.96 234.36 280.76 ;
      RECT 233.78 283.36 234.36 284.16 ;
      RECT 233.78 286.76 234.36 287.56 ;
      RECT 233.78 290.16 234.36 290.96 ;
      RECT 233.78 293.56 234.36 294.36 ;
      RECT 233.78 296.96 234.36 297.76 ;
      RECT 233.78 300.36 234.36 301.16 ;
      RECT 233.78 303.76 234.36 304.56 ;
      RECT 233.78 307.16 234.36 307.96 ;
      RECT 233.78 310.56 234.36 311.36 ;
      RECT 233.78 313.96 234.36 314.76 ;
      RECT 233.78 317.36 234.36 318.16 ;
      RECT 233.78 320.76 234.36 321.56 ;
      RECT 233.78 324.16 234.36 324.96 ;
      RECT 233.78 327.56 234.36 328.36 ;
      RECT 233.78 330.96 234.36 331.76 ;
      RECT 233.78 334.36 234.36 335.16 ;
      RECT 233.78 337.76 234.36 338.56 ;
      RECT 233.78 341.16 234.36 341.96 ;
      RECT 233.78 344.56 234.36 345.36 ;
      RECT 233.78 347.96 234.36 348.76 ;
      RECT 233.78 351.36 234.36 352.16 ;
      RECT 233.78 354.76 234.36 355.56 ;
      RECT 233.78 358.16 234.36 358.96 ;
      RECT 233.78 361.56 234.36 362.36 ;
      RECT 233.78 364.96 234.36 365.76 ;
      RECT 233.78 368.36 234.36 369.16 ;
      RECT 233.78 371.76 234.36 372.56 ;
      RECT 233.78 375.16 234.36 375.96 ;
      RECT 233.78 378.56 234.36 379.36 ;
      RECT 233.78 381.96 234.36 382.76 ;
      RECT 233.78 385.36 234.36 386.16 ;
      RECT 233.78 388.76 234.36 389.56 ;
      RECT 233.78 392.16 234.36 392.96 ;
      RECT 233.78 395.56 234.36 396.36 ;
      RECT 233.78 398.96 234.36 399.76 ;
      RECT 233.78 402.36 234.36 403.16 ;
      RECT 233.78 405.76 234.36 406.56 ;
      RECT 233.78 409.16 234.36 409.96 ;
      RECT 233.78 412.56 234.36 413.36 ;
      RECT 233.78 415.96 234.36 416.76 ;
      RECT 233.78 419.36 234.36 420.16 ;
      RECT 233.78 422.76 234.36 423.56 ;
      RECT 233.78 426.16 234.36 426.96 ;
      RECT 233.78 429.56 234.36 430.36 ;
      RECT 233.78 432.96 234.36 433.76 ;
      RECT 233.78 436.36 234.36 437.16 ;
      RECT 233.78 439.76 234.36 440.56 ;
      RECT 233.78 443.16 234.36 443.96 ;
      RECT 233.78 446.56 234.36 447.36 ;
      RECT 233.78 449.96 234.36 450.76 ;
      RECT 233.78 453.36 234.36 454.16 ;
      RECT 233.78 456.76 234.36 457.56 ;
      RECT 233.78 460.16 234.36 460.96 ;
      RECT 233.78 463.56 234.36 464.36 ;
      RECT 233.78 466.96 234.36 467.76 ;
      RECT 233.78 470.36 234.36 471.16 ;
      RECT 233.78 473.76 234.36 474.56 ;
      RECT 233.78 477.16 234.36 477.96 ;
      RECT 233.78 480.56 234.36 481.36 ;
      RECT 233.78 483.96 234.36 484.76 ;
      RECT 233.78 487.36 234.36 488.16 ;
      RECT 233.78 490.76 234.36 491.56 ;
      RECT 233.78 494.16 234.36 494.96 ;
      RECT 233.78 497.56 234.36 498.36 ;
      RECT 233.78 500.96 234.36 501.76 ;
      RECT 233.78 504.36 234.36 505.16 ;
      RECT 233.78 505.6 234.36 506 ;
      RECT 233.78 509 234.36 509.8 ;
      RECT 233.6 9.34 233.85 9.78 ;
      RECT 233.57 10.92 233.85 11.4 ;
      RECT 233.58 14.87 233.85 15.29 ;
      RECT 233.57 18.87 233.85 19.35 ;
      RECT 231.19 6.24 233.19 6.84 ;
      RECT 232.09 36.22 232.29 36.95 ;
      RECT 232.11 29.32 232.27 34.08 ;
      RECT 232.11 39.34 232.27 46.59 ;
      RECT 232.11 47.59 232.27 51.92 ;
      RECT 232.11 52.64 232.27 56.5 ;
      RECT 231.79 47.88 231.95 51.16 ;
      RECT 231.63 57.79 231.79 62.72 ;
      RECT 231.39 29.97 231.55 32.28 ;
      RECT 231.39 35.23 231.55 36.31 ;
      RECT 231.39 37.11 231.55 38.19 ;
      RECT 231.39 41.14 231.55 43.45 ;
      RECT 223.47 15.46 231.31 16.9 ;
      RECT 231.15 57.79 231.31 62.72 ;
      RECT 230.79 56.99 231.19 57.29 ;
      RECT 230.91 29.97 231.07 34.08 ;
      RECT 230.91 39.34 231.07 43.45 ;
      RECT 230.83 48.24 230.99 50.5 ;
      RECT 230.67 57.79 230.83 67.9 ;
      RECT 228.81 6.24 230.79 6.84 ;
      RECT 228.79 510.54 230.79 510.94 ;
      RECT 230.43 29.97 230.59 32.28 ;
      RECT 230.43 35.23 230.59 36.31 ;
      RECT 230.43 37.11 230.59 38.19 ;
      RECT 230.43 41.14 230.59 43.45 ;
      RECT 224.37 21.67 230.41 21.95 ;
      RECT 229.69 36.21 229.89 36.95 ;
      RECT 229.71 29.32 229.87 34.08 ;
      RECT 229.71 39.34 229.87 46.59 ;
      RECT 229.71 47.59 229.87 51.11 ;
      RECT 229.71 51.34 229.87 53.67 ;
      RECT 229.71 54.16 229.87 56.5 ;
      RECT 228.99 29.97 229.15 32.28 ;
      RECT 228.99 35.23 229.15 36.31 ;
      RECT 228.99 37.11 229.15 38.19 ;
      RECT 228.99 41.14 229.15 43.45 ;
      RECT 228.75 57.79 228.91 67.9 ;
      RECT 228.39 56.99 228.79 57.29 ;
      RECT 228.59 48.24 228.75 50.5 ;
      RECT 228.51 29.97 228.67 34.08 ;
      RECT 228.51 39.34 228.67 43.45 ;
      RECT 228.27 57.79 228.43 62.72 ;
      RECT 226.41 6.24 228.39 6.84 ;
      RECT 228.03 29.97 228.19 32.28 ;
      RECT 228.03 35.23 228.19 36.31 ;
      RECT 228.03 37.11 228.19 38.19 ;
      RECT 228.03 41.14 228.19 43.45 ;
      RECT 227.79 57.79 227.95 62.72 ;
      RECT 227.63 47.88 227.79 51.16 ;
      RECT 227.11 9.36 227.67 9.52 ;
      RECT 227.11 11.3 227.67 11.46 ;
      RECT 227.11 14.68 227.67 14.84 ;
      RECT 227.11 19.63 227.67 19.79 ;
      RECT 227.29 36.21 227.49 36.95 ;
      RECT 227.31 29.32 227.47 34.08 ;
      RECT 227.31 39.34 227.47 46.59 ;
      RECT 227.31 47.59 227.47 51.92 ;
      RECT 227.31 52.64 227.47 56.5 ;
      RECT 226.99 47.88 227.15 51.16 ;
      RECT 226.83 57.79 226.99 62.72 ;
      RECT 226.59 29.97 226.75 32.28 ;
      RECT 226.59 35.23 226.75 36.31 ;
      RECT 226.59 37.11 226.75 38.19 ;
      RECT 226.59 41.14 226.75 43.45 ;
      RECT 226.35 57.79 226.51 62.72 ;
      RECT 225.99 56.99 226.39 57.29 ;
      RECT 226.11 29.97 226.27 34.08 ;
      RECT 226.11 39.34 226.27 43.45 ;
      RECT 226.03 48.24 226.19 50.5 ;
      RECT 225.87 57.79 226.03 67.9 ;
      RECT 224.01 6.24 225.99 6.84 ;
      RECT 223.99 510.54 225.99 510.94 ;
      RECT 225.63 29.97 225.79 32.28 ;
      RECT 225.63 35.23 225.79 36.31 ;
      RECT 225.63 37.11 225.79 38.19 ;
      RECT 225.63 41.14 225.79 43.45 ;
      RECT 224.89 36.21 225.09 36.95 ;
      RECT 224.91 29.32 225.07 34.08 ;
      RECT 224.91 39.34 225.07 46.59 ;
      RECT 224.91 47.59 225.07 51.11 ;
      RECT 224.91 51.34 225.07 53.67 ;
      RECT 224.91 54.16 225.07 56.5 ;
      RECT 224.19 29.97 224.35 32.28 ;
      RECT 224.19 35.23 224.35 36.31 ;
      RECT 224.19 37.11 224.35 38.19 ;
      RECT 224.19 41.14 224.35 43.45 ;
      RECT 223.95 57.79 224.11 67.9 ;
      RECT 223.59 56.99 223.99 57.29 ;
      RECT 223.79 48.24 223.95 50.5 ;
      RECT 223.71 29.97 223.87 34.08 ;
      RECT 223.71 39.34 223.87 43.45 ;
      RECT 223.47 57.79 223.63 62.72 ;
      RECT 221.59 6.24 223.59 6.84 ;
      RECT 223.23 29.97 223.39 32.28 ;
      RECT 223.23 35.23 223.39 36.31 ;
      RECT 223.23 37.11 223.39 38.19 ;
      RECT 223.23 41.14 223.39 43.45 ;
      RECT 222.99 57.79 223.15 62.72 ;
      RECT 222.83 47.88 222.99 51.16 ;
      RECT 222.49 36.21 222.69 36.95 ;
      RECT 222.51 21.45 222.67 24.52 ;
      RECT 222.51 29.32 222.67 34.08 ;
      RECT 222.51 39.34 222.67 46.59 ;
      RECT 222.51 47.59 222.67 51.92 ;
      RECT 222.51 52.64 222.67 56.5 ;
      RECT 221.84 8.96 222.35 9.17 ;
      RECT 222.19 47.83 222.35 51.16 ;
      RECT 222.05 15.09 222.33 15.41 ;
      RECT 222.03 57.79 222.19 62.72 ;
      RECT 221.83 12.28 222.15 12.76 ;
      RECT 221.87 21.73 222.03 22.33 ;
      RECT 221.87 22.49 222.03 23.06 ;
      RECT 221.79 29.97 221.95 32.28 ;
      RECT 221.79 35.23 221.95 36.31 ;
      RECT 221.79 37.11 221.95 38.19 ;
      RECT 221.79 41.14 221.95 43.45 ;
      RECT 221.55 57.79 221.71 62.72 ;
      RECT 221.19 56.99 221.59 57.29 ;
      RECT 220.41 13.4 221.53 13.56 ;
      RECT 221.31 29.97 221.47 34.08 ;
      RECT 221.31 39.34 221.47 43.45 ;
      RECT 221.3 26.68 221.46 28.17 ;
      RECT 221.23 48.24 221.39 50.5 ;
      RECT 221.03 10.76 221.35 11.16 ;
      RECT 220.61 10 221.33 10.18 ;
      RECT 221.07 57.79 221.23 67.9 ;
      RECT 219.21 6.24 221.19 6.84 ;
      RECT 219.19 510.54 221.19 510.94 ;
      RECT 220.83 29.97 220.99 32.28 ;
      RECT 220.83 35.23 220.99 36.31 ;
      RECT 220.83 37.11 220.99 38.19 ;
      RECT 220.83 41.14 220.99 43.45 ;
      RECT 220.52 17 220.68 18.12 ;
      RECT 220.09 36.21 220.29 36.95 ;
      RECT 220.11 29.32 220.27 34.08 ;
      RECT 220.11 39.34 220.27 46.59 ;
      RECT 220.11 47.59 220.27 51.11 ;
      RECT 220.11 51.34 220.27 53.67 ;
      RECT 220.11 54.16 220.27 56.5 ;
      RECT 219.79 23.54 220.23 23.81 ;
      RECT 219.88 15.33 220.04 15.89 ;
      RECT 219.32 28.33 219.88 28.49 ;
      RECT 219.39 25.51 219.63 26.2 ;
      RECT 219.39 29.97 219.55 32.28 ;
      RECT 219.39 35.23 219.55 36.31 ;
      RECT 219.39 37.11 219.55 38.19 ;
      RECT 219.39 41.14 219.55 43.45 ;
      RECT 219.15 57.79 219.31 67.9 ;
      RECT 218.79 56.99 219.19 57.29 ;
      RECT 219 16.21 219.16 18.62 ;
      RECT 218.99 48.24 219.15 50.5 ;
      RECT 218.91 29.97 219.07 34.08 ;
      RECT 218.91 39.34 219.07 43.45 ;
      RECT 218.85 14.84 219.01 16.05 ;
      RECT 218.67 57.79 218.83 62.72 ;
      RECT 217.29 6.24 218.79 6.84 ;
      RECT 218.43 29.97 218.59 32.28 ;
      RECT 218.43 35.23 218.59 36.31 ;
      RECT 218.43 37.11 218.59 38.19 ;
      RECT 218.43 41.14 218.59 43.45 ;
      RECT 218.19 57.79 218.35 62.72 ;
      RECT 217.97 19.63 218.29 20.04 ;
      RECT 218.03 47.88 218.19 51.16 ;
      RECT 217.53 13.8 218.09 13.96 ;
      RECT 217.41 13.32 217.89 13.56 ;
      RECT 217.69 36.21 217.89 36.95 ;
      RECT 217.71 26.38 217.87 27.85 ;
      RECT 217.71 29.32 217.87 34.08 ;
      RECT 217.71 39.34 217.87 46.59 ;
      RECT 217.71 47.59 217.87 51.92 ;
      RECT 217.71 52.64 217.87 56.5 ;
      RECT 217.39 47.88 217.55 51.16 ;
      RECT 216.99 16.47 217.41 17.1 ;
      RECT 217.23 57.79 217.39 62.72 ;
      RECT 216.99 29.97 217.15 32.28 ;
      RECT 216.99 35.23 217.15 36.31 ;
      RECT 216.99 37.11 217.15 38.19 ;
      RECT 216.99 41.14 217.15 43.45 ;
      RECT 216.75 57.79 216.91 62.72 ;
      RECT 216.39 56.99 216.79 57.29 ;
      RECT 216.51 29.97 216.67 34.08 ;
      RECT 216.51 39.34 216.67 43.45 ;
      RECT 216.43 48.24 216.59 50.5 ;
      RECT 216.27 57.79 216.43 67.9 ;
      RECT 214.39 510.54 216.39 510.94 ;
      RECT 215.7 28.33 216.26 28.49 ;
      RECT 215.95 25.51 216.19 26.2 ;
      RECT 216.03 29.97 216.19 32.28 ;
      RECT 216.03 35.23 216.19 36.31 ;
      RECT 216.03 37.11 216.19 38.19 ;
      RECT 216.03 41.14 216.19 43.45 ;
      RECT 214.89 6.24 215.89 6.84 ;
      RECT 215.35 23.54 215.79 23.81 ;
      RECT 215.29 36.21 215.49 36.95 ;
      RECT 215.31 29.32 215.47 34.08 ;
      RECT 215.31 39.34 215.47 46.59 ;
      RECT 215.31 47.59 215.47 51.11 ;
      RECT 215.31 51.34 215.47 53.67 ;
      RECT 215.31 54.16 215.47 56.5 ;
      RECT 215.11 21.85 215.27 22.91 ;
      RECT 215.08 7.58 215.24 8.64 ;
      RECT 215.04 20.65 215.2 21.69 ;
      RECT 213.73 16.8 214.75 17.08 ;
      RECT 214.59 29.97 214.75 32.28 ;
      RECT 214.59 35.23 214.75 36.31 ;
      RECT 214.59 37.11 214.75 38.19 ;
      RECT 214.59 41.14 214.75 43.45 ;
      RECT 214.27 15.32 214.67 15.64 ;
      RECT 214.35 57.79 214.51 67.9 ;
      RECT 213.99 56.99 214.39 57.29 ;
      RECT 214.2 8.04 214.36 8.6 ;
      RECT 214.19 48.24 214.35 50.5 ;
      RECT 213.73 16.12 214.29 16.28 ;
      RECT 214.12 26.68 214.28 28.17 ;
      RECT 214.11 29.97 214.27 34.08 ;
      RECT 214.11 39.34 214.27 43.45 ;
      RECT 213.87 11.52 214.03 13.07 ;
      RECT 213.87 57.79 214.03 62.72 ;
      RECT 213.63 29.97 213.79 32.28 ;
      RECT 213.63 35.23 213.79 36.31 ;
      RECT 213.63 37.11 213.79 38.19 ;
      RECT 213.63 41.14 213.79 43.45 ;
      RECT 213.51 13.11 213.67 13.67 ;
      RECT 213.39 57.79 213.55 62.72 ;
      RECT 212.59 6.24 213.39 6.84 ;
      RECT 213.23 47.88 213.39 51.16 ;
      RECT 212.89 36.21 213.09 36.95 ;
      RECT 212.91 21.45 213.07 24.52 ;
      RECT 212.91 29.32 213.07 34.08 ;
      RECT 212.91 39.34 213.07 46.59 ;
      RECT 212.91 47.59 213.07 51.92 ;
      RECT 212.91 52.64 213.07 56.5 ;
      RECT 212.59 47.88 212.75 51.16 ;
      RECT 212.43 57.79 212.59 62.72 ;
      RECT 212.31 13.11 212.47 13.67 ;
      RECT 212.19 29.97 212.35 32.28 ;
      RECT 212.19 35.23 212.35 36.31 ;
      RECT 212.19 37.11 212.35 38.19 ;
      RECT 212.19 41.14 212.35 43.45 ;
      RECT 211.69 16.12 212.25 16.28 ;
      RECT 211.23 16.8 212.25 17.08 ;
      RECT 211.95 11.52 212.11 13.07 ;
      RECT 211.95 57.79 212.11 62.72 ;
      RECT 211.59 56.99 211.99 57.29 ;
      RECT 211.71 29.97 211.87 34.08 ;
      RECT 211.71 39.34 211.87 43.45 ;
      RECT 211.7 26.68 211.86 28.17 ;
      RECT 211.63 48.24 211.79 50.5 ;
      RECT 211.62 8.04 211.78 8.6 ;
      RECT 211.31 15.32 211.71 15.64 ;
      RECT 211.47 57.79 211.63 67.9 ;
      RECT 209.59 510.54 211.59 510.94 ;
      RECT 211.23 29.97 211.39 32.28 ;
      RECT 211.23 35.23 211.39 36.31 ;
      RECT 211.23 37.11 211.39 38.19 ;
      RECT 211.23 41.14 211.39 43.45 ;
      RECT 210.09 6.24 211.09 6.84 ;
      RECT 210.78 20.65 210.94 21.69 ;
      RECT 210.74 7.58 210.9 8.64 ;
      RECT 210.71 21.85 210.87 22.91 ;
      RECT 210.49 36.21 210.69 36.95 ;
      RECT 210.51 29.32 210.67 34.08 ;
      RECT 210.51 39.34 210.67 46.59 ;
      RECT 210.51 47.59 210.67 51.11 ;
      RECT 210.51 51.34 210.67 53.67 ;
      RECT 210.51 54.16 210.67 56.5 ;
      RECT 210.19 23.54 210.63 23.81 ;
      RECT 209.72 28.33 210.28 28.49 ;
      RECT 209.79 25.51 210.03 26.2 ;
      RECT 209.79 29.97 209.95 32.28 ;
      RECT 209.79 35.23 209.95 36.31 ;
      RECT 209.79 37.11 209.95 38.19 ;
      RECT 209.79 41.14 209.95 43.45 ;
      RECT 209.55 57.79 209.71 67.9 ;
      RECT 209.19 56.99 209.59 57.29 ;
      RECT 209.39 48.24 209.55 50.5 ;
      RECT 209.31 29.97 209.47 34.08 ;
      RECT 209.31 39.34 209.47 43.45 ;
      RECT 209.07 57.79 209.23 62.72 ;
      RECT 208.57 16.47 208.99 17.1 ;
      RECT 208.83 29.97 208.99 32.28 ;
      RECT 208.83 35.23 208.99 36.31 ;
      RECT 208.83 37.11 208.99 38.19 ;
      RECT 208.83 41.14 208.99 43.45 ;
      RECT 208.59 57.79 208.75 62.72 ;
      RECT 207.19 6.24 208.69 6.84 ;
      RECT 208.43 47.88 208.59 51.16 ;
      RECT 208.09 13.32 208.57 13.56 ;
      RECT 207.89 13.8 208.45 13.96 ;
      RECT 208.09 36.21 208.29 36.95 ;
      RECT 208.11 26.38 208.27 27.85 ;
      RECT 208.11 29.32 208.27 34.08 ;
      RECT 208.11 39.34 208.27 46.59 ;
      RECT 208.11 47.59 208.27 51.92 ;
      RECT 208.11 52.64 208.27 56.5 ;
      RECT 207.69 19.63 208.01 20.04 ;
      RECT 207.79 47.88 207.95 51.16 ;
      RECT 207.63 57.79 207.79 62.72 ;
      RECT 207.39 29.97 207.55 32.28 ;
      RECT 207.39 35.23 207.55 36.31 ;
      RECT 207.39 37.11 207.55 38.19 ;
      RECT 207.39 41.14 207.55 43.45 ;
      RECT 207.15 57.79 207.31 62.72 ;
      RECT 206.79 56.99 207.19 57.29 ;
      RECT 206.97 14.84 207.13 16.05 ;
      RECT 206.91 29.97 207.07 34.08 ;
      RECT 206.91 39.34 207.07 43.45 ;
      RECT 206.83 48.24 206.99 50.5 ;
      RECT 206.82 16.21 206.98 18.62 ;
      RECT 206.67 57.79 206.83 67.9 ;
      RECT 204.79 510.54 206.79 510.94 ;
      RECT 204.79 6.24 206.76 6.84 ;
      RECT 206.1 28.33 206.66 28.49 ;
      RECT 206.35 25.51 206.59 26.2 ;
      RECT 206.43 29.97 206.59 32.28 ;
      RECT 206.43 35.23 206.59 36.31 ;
      RECT 206.43 37.11 206.59 38.19 ;
      RECT 206.43 41.14 206.59 43.45 ;
      RECT 205.75 23.54 206.19 23.81 ;
      RECT 205.94 15.33 206.1 15.89 ;
      RECT 205.69 36.21 205.89 36.95 ;
      RECT 205.71 29.32 205.87 34.08 ;
      RECT 205.71 39.34 205.87 46.59 ;
      RECT 205.71 47.59 205.87 51.11 ;
      RECT 205.71 51.34 205.87 53.67 ;
      RECT 205.71 54.16 205.87 56.5 ;
      RECT 204.45 13.4 205.57 13.56 ;
      RECT 205.3 17 205.46 18.12 ;
      RECT 204.65 10 205.37 10.18 ;
      RECT 204.99 29.97 205.15 32.28 ;
      RECT 204.99 35.23 205.15 36.31 ;
      RECT 204.99 37.11 205.15 38.19 ;
      RECT 204.99 41.14 205.15 43.45 ;
      RECT 204.63 10.76 204.95 11.16 ;
      RECT 204.75 57.79 204.91 67.9 ;
      RECT 204.39 56.99 204.79 57.29 ;
      RECT 204.59 48.24 204.75 50.5 ;
      RECT 204.52 26.68 204.68 28.17 ;
      RECT 204.51 29.97 204.67 34.08 ;
      RECT 204.51 39.34 204.67 43.45 ;
      RECT 204.27 57.79 204.43 62.72 ;
      RECT 202.39 6.24 204.39 6.84 ;
      RECT 204.03 29.97 204.19 32.28 ;
      RECT 204.03 35.23 204.19 36.31 ;
      RECT 204.03 37.11 204.19 38.19 ;
      RECT 204.03 41.14 204.19 43.45 ;
      RECT 203.83 12.28 204.15 12.76 ;
      RECT 203.63 8.96 204.14 9.17 ;
      RECT 203.95 21.73 204.11 22.33 ;
      RECT 203.95 22.49 204.11 23.06 ;
      RECT 203.79 57.79 203.95 62.72 ;
      RECT 203.65 15.09 203.93 15.41 ;
      RECT 203.63 47.88 203.79 51.16 ;
      RECT 203.29 36.21 203.49 36.95 ;
      RECT 203.31 21.45 203.47 24.52 ;
      RECT 203.31 29.32 203.47 34.08 ;
      RECT 203.31 39.34 203.47 46.59 ;
      RECT 203.31 47.59 203.47 51.92 ;
      RECT 203.31 52.64 203.47 56.5 ;
      RECT 202.99 47.83 203.15 51.16 ;
      RECT 202.83 57.79 202.99 62.72 ;
      RECT 202.59 29.97 202.75 32.28 ;
      RECT 202.59 35.23 202.75 36.31 ;
      RECT 202.59 37.11 202.75 38.19 ;
      RECT 202.59 41.14 202.75 43.45 ;
      RECT 194.67 15.46 202.51 16.9 ;
      RECT 202.35 57.79 202.51 62.72 ;
      RECT 201.99 56.99 202.39 57.29 ;
      RECT 202.11 29.97 202.27 34.08 ;
      RECT 202.11 39.34 202.27 43.45 ;
      RECT 202.03 48.24 202.19 50.5 ;
      RECT 201.87 57.79 202.03 67.9 ;
      RECT 199.99 510.54 201.99 510.94 ;
      RECT 199.99 6.24 201.97 6.84 ;
      RECT 201.63 29.97 201.79 32.28 ;
      RECT 201.63 35.23 201.79 36.31 ;
      RECT 201.63 37.11 201.79 38.19 ;
      RECT 201.63 41.14 201.79 43.45 ;
      RECT 195.57 21.67 201.61 21.95 ;
      RECT 200.89 36.21 201.09 36.95 ;
      RECT 200.91 29.32 201.07 34.08 ;
      RECT 200.91 39.34 201.07 46.59 ;
      RECT 200.91 47.59 201.07 51.11 ;
      RECT 200.91 51.34 201.07 53.67 ;
      RECT 200.91 54.16 201.07 56.5 ;
      RECT 200.19 29.97 200.35 32.28 ;
      RECT 200.19 35.23 200.35 36.31 ;
      RECT 200.19 37.11 200.35 38.19 ;
      RECT 200.19 41.14 200.35 43.45 ;
      RECT 199.95 57.79 200.11 67.9 ;
      RECT 199.59 56.99 199.99 57.29 ;
      RECT 199.79 48.24 199.95 50.5 ;
      RECT 199.71 29.97 199.87 34.08 ;
      RECT 199.71 39.34 199.87 43.45 ;
      RECT 199.47 57.79 199.63 62.72 ;
      RECT 197.59 6.24 199.57 6.84 ;
      RECT 199.23 29.97 199.39 32.28 ;
      RECT 199.23 35.23 199.39 36.31 ;
      RECT 199.23 37.11 199.39 38.19 ;
      RECT 199.23 41.14 199.39 43.45 ;
      RECT 198.99 57.79 199.15 62.72 ;
      RECT 198.83 47.88 198.99 51.16 ;
      RECT 198.31 9.36 198.87 9.52 ;
      RECT 198.31 11.3 198.87 11.46 ;
      RECT 198.31 14.68 198.87 14.84 ;
      RECT 198.31 19.63 198.87 19.79 ;
      RECT 198.49 36.21 198.69 36.95 ;
      RECT 198.51 29.32 198.67 34.08 ;
      RECT 198.51 39.34 198.67 46.59 ;
      RECT 198.51 47.59 198.67 51.92 ;
      RECT 198.51 52.64 198.67 56.5 ;
      RECT 198.19 47.88 198.35 51.16 ;
      RECT 198.03 57.79 198.19 62.72 ;
      RECT 197.79 29.97 197.95 32.28 ;
      RECT 197.79 35.23 197.95 36.31 ;
      RECT 197.79 37.11 197.95 38.19 ;
      RECT 197.79 41.14 197.95 43.45 ;
      RECT 197.55 57.79 197.71 62.72 ;
      RECT 197.19 56.99 197.59 57.29 ;
      RECT 197.31 29.97 197.47 34.08 ;
      RECT 197.31 39.34 197.47 43.45 ;
      RECT 197.23 48.24 197.39 50.5 ;
      RECT 197.07 57.79 197.23 67.9 ;
      RECT 195.19 510.54 197.19 510.94 ;
      RECT 195.19 6.24 197.17 6.84 ;
      RECT 196.83 29.97 196.99 32.28 ;
      RECT 196.83 35.23 196.99 36.31 ;
      RECT 196.83 37.11 196.99 38.19 ;
      RECT 196.83 41.14 196.99 43.45 ;
      RECT 196.09 36.21 196.29 36.95 ;
      RECT 196.11 29.32 196.27 34.08 ;
      RECT 196.11 39.34 196.27 46.59 ;
      RECT 196.11 47.59 196.27 51.11 ;
      RECT 196.11 51.34 196.27 53.67 ;
      RECT 196.11 54.16 196.27 56.5 ;
      RECT 195.39 29.97 195.55 32.28 ;
      RECT 195.39 35.23 195.55 36.31 ;
      RECT 195.39 37.11 195.55 38.19 ;
      RECT 195.39 41.14 195.55 43.45 ;
      RECT 195.15 57.79 195.31 67.9 ;
      RECT 194.79 56.99 195.19 57.29 ;
      RECT 194.99 48.24 195.15 50.5 ;
      RECT 194.91 29.97 195.07 34.08 ;
      RECT 194.91 39.34 195.07 43.45 ;
      RECT 194.67 57.79 194.83 62.72 ;
      RECT 194.43 29.97 194.59 32.28 ;
      RECT 194.43 35.23 194.59 36.31 ;
      RECT 194.43 37.11 194.59 38.19 ;
      RECT 194.43 41.14 194.59 43.45 ;
      RECT 194.19 57.79 194.35 62.72 ;
      RECT 194.03 47.88 194.19 51.16 ;
      RECT 193.69 36.21 193.89 36.95 ;
      RECT 193.71 29.32 193.87 34.08 ;
      RECT 193.71 39.34 193.87 46.59 ;
      RECT 193.71 47.59 193.87 51.92 ;
      RECT 193.71 52.64 193.87 56.5 ;
      RECT 193.09 36.11 193.29 58.16 ;
      RECT 193.11 8.48 193.27 10.44 ;
      RECT 193.11 17.36 193.27 17.92 ;
      RECT 193.11 20.74 193.27 27.31 ;
      RECT 192.49 36.22 192.69 36.95 ;
      RECT 192.51 29.32 192.67 34.08 ;
      RECT 192.51 39.34 192.67 46.59 ;
      RECT 192.51 47.59 192.67 51.92 ;
      RECT 192.51 52.64 192.67 56.5 ;
      RECT 192.19 47.88 192.35 51.16 ;
      RECT 192.03 57.79 192.19 62.72 ;
      RECT 191.79 29.97 191.95 32.28 ;
      RECT 191.79 35.23 191.95 36.31 ;
      RECT 191.79 37.11 191.95 38.19 ;
      RECT 191.79 41.14 191.95 43.45 ;
      RECT 183.87 15.46 191.71 16.9 ;
      RECT 191.55 57.79 191.71 62.72 ;
      RECT 191.19 56.99 191.59 57.29 ;
      RECT 191.31 29.97 191.47 34.08 ;
      RECT 191.31 39.34 191.47 43.45 ;
      RECT 191.23 48.24 191.39 50.5 ;
      RECT 191.07 57.79 191.23 67.9 ;
      RECT 189.21 6.24 191.19 6.84 ;
      RECT 189.19 510.54 191.19 510.94 ;
      RECT 190.83 29.97 190.99 32.28 ;
      RECT 190.83 35.23 190.99 36.31 ;
      RECT 190.83 37.11 190.99 38.19 ;
      RECT 190.83 41.14 190.99 43.45 ;
      RECT 184.77 21.67 190.81 21.95 ;
      RECT 190.09 36.21 190.29 36.95 ;
      RECT 190.11 29.32 190.27 34.08 ;
      RECT 190.11 39.34 190.27 46.59 ;
      RECT 190.11 47.59 190.27 51.11 ;
      RECT 190.11 51.34 190.27 53.67 ;
      RECT 190.11 54.16 190.27 56.5 ;
      RECT 189.39 29.97 189.55 32.28 ;
      RECT 189.39 35.23 189.55 36.31 ;
      RECT 189.39 37.11 189.55 38.19 ;
      RECT 189.39 41.14 189.55 43.45 ;
      RECT 189.15 57.79 189.31 67.9 ;
      RECT 188.79 56.99 189.19 57.29 ;
      RECT 188.99 48.24 189.15 50.5 ;
      RECT 188.91 29.97 189.07 34.08 ;
      RECT 188.91 39.34 189.07 43.45 ;
      RECT 188.67 57.79 188.83 62.72 ;
      RECT 186.81 6.24 188.79 6.84 ;
      RECT 188.43 29.97 188.59 32.28 ;
      RECT 188.43 35.23 188.59 36.31 ;
      RECT 188.43 37.11 188.59 38.19 ;
      RECT 188.43 41.14 188.59 43.45 ;
      RECT 188.19 57.79 188.35 62.72 ;
      RECT 188.03 47.88 188.19 51.16 ;
      RECT 187.51 9.36 188.07 9.52 ;
      RECT 187.51 11.3 188.07 11.46 ;
      RECT 187.51 14.68 188.07 14.84 ;
      RECT 187.51 19.63 188.07 19.79 ;
      RECT 187.69 36.21 187.89 36.95 ;
      RECT 187.71 29.32 187.87 34.08 ;
      RECT 187.71 39.34 187.87 46.59 ;
      RECT 187.71 47.59 187.87 51.92 ;
      RECT 187.71 52.64 187.87 56.5 ;
      RECT 187.39 47.88 187.55 51.16 ;
      RECT 187.23 57.79 187.39 62.72 ;
      RECT 186.99 29.97 187.15 32.28 ;
      RECT 186.99 35.23 187.15 36.31 ;
      RECT 186.99 37.11 187.15 38.19 ;
      RECT 186.99 41.14 187.15 43.45 ;
      RECT 186.75 57.79 186.91 62.72 ;
      RECT 186.39 56.99 186.79 57.29 ;
      RECT 186.51 29.97 186.67 34.08 ;
      RECT 186.51 39.34 186.67 43.45 ;
      RECT 186.43 48.24 186.59 50.5 ;
      RECT 186.27 57.79 186.43 67.9 ;
      RECT 184.41 6.24 186.39 6.84 ;
      RECT 184.39 510.54 186.39 510.94 ;
      RECT 186.03 29.97 186.19 32.28 ;
      RECT 186.03 35.23 186.19 36.31 ;
      RECT 186.03 37.11 186.19 38.19 ;
      RECT 186.03 41.14 186.19 43.45 ;
      RECT 185.29 36.21 185.49 36.95 ;
      RECT 185.31 29.32 185.47 34.08 ;
      RECT 185.31 39.34 185.47 46.59 ;
      RECT 185.31 47.59 185.47 51.11 ;
      RECT 185.31 51.34 185.47 53.67 ;
      RECT 185.31 54.16 185.47 56.5 ;
      RECT 184.59 29.97 184.75 32.28 ;
      RECT 184.59 35.23 184.75 36.31 ;
      RECT 184.59 37.11 184.75 38.19 ;
      RECT 184.59 41.14 184.75 43.45 ;
      RECT 184.35 57.79 184.51 67.9 ;
      RECT 183.99 56.99 184.39 57.29 ;
      RECT 184.19 48.24 184.35 50.5 ;
      RECT 184.11 29.97 184.27 34.08 ;
      RECT 184.11 39.34 184.27 43.45 ;
      RECT 183.87 57.79 184.03 62.72 ;
      RECT 181.99 6.24 183.99 6.84 ;
      RECT 183.63 29.97 183.79 32.28 ;
      RECT 183.63 35.23 183.79 36.31 ;
      RECT 183.63 37.11 183.79 38.19 ;
      RECT 183.63 41.14 183.79 43.45 ;
      RECT 183.39 57.79 183.55 62.72 ;
      RECT 183.23 47.88 183.39 51.16 ;
      RECT 182.89 36.21 183.09 36.95 ;
      RECT 182.91 21.45 183.07 24.52 ;
      RECT 182.91 29.32 183.07 34.08 ;
      RECT 182.91 39.34 183.07 46.59 ;
      RECT 182.91 47.59 183.07 51.92 ;
      RECT 182.91 52.64 183.07 56.5 ;
      RECT 182.24 8.96 182.75 9.17 ;
      RECT 182.59 47.83 182.75 51.16 ;
      RECT 182.45 15.09 182.73 15.41 ;
      RECT 182.43 57.79 182.59 62.72 ;
      RECT 182.23 12.28 182.55 12.76 ;
      RECT 182.27 21.73 182.43 22.33 ;
      RECT 182.27 22.49 182.43 23.06 ;
      RECT 182.19 29.97 182.35 32.28 ;
      RECT 182.19 35.23 182.35 36.31 ;
      RECT 182.19 37.11 182.35 38.19 ;
      RECT 182.19 41.14 182.35 43.45 ;
      RECT 181.95 57.79 182.11 62.72 ;
      RECT 181.59 56.99 181.99 57.29 ;
      RECT 180.81 13.4 181.93 13.56 ;
      RECT 181.71 29.97 181.87 34.08 ;
      RECT 181.71 39.34 181.87 43.45 ;
      RECT 181.7 26.68 181.86 28.17 ;
      RECT 181.63 48.24 181.79 50.5 ;
      RECT 181.43 10.76 181.75 11.16 ;
      RECT 181.01 10 181.73 10.18 ;
      RECT 181.47 57.79 181.63 67.9 ;
      RECT 179.62 6.24 181.59 6.84 ;
      RECT 179.59 510.54 181.59 510.94 ;
      RECT 181.23 29.97 181.39 32.28 ;
      RECT 181.23 35.23 181.39 36.31 ;
      RECT 181.23 37.11 181.39 38.19 ;
      RECT 181.23 41.14 181.39 43.45 ;
      RECT 180.92 17 181.08 18.12 ;
      RECT 180.49 36.21 180.69 36.95 ;
      RECT 180.51 29.32 180.67 34.08 ;
      RECT 180.51 39.34 180.67 46.59 ;
      RECT 180.51 47.59 180.67 51.11 ;
      RECT 180.51 51.34 180.67 53.67 ;
      RECT 180.51 54.16 180.67 56.5 ;
      RECT 180.19 23.54 180.63 23.81 ;
      RECT 180.28 15.33 180.44 15.89 ;
      RECT 179.72 28.33 180.28 28.49 ;
      RECT 179.79 25.51 180.03 26.2 ;
      RECT 179.79 29.97 179.95 32.28 ;
      RECT 179.79 35.23 179.95 36.31 ;
      RECT 179.79 37.11 179.95 38.19 ;
      RECT 179.79 41.14 179.95 43.45 ;
      RECT 179.55 57.79 179.71 67.9 ;
      RECT 179.19 56.99 179.59 57.29 ;
      RECT 179.4 16.21 179.56 18.62 ;
      RECT 179.39 48.24 179.55 50.5 ;
      RECT 179.31 29.97 179.47 34.08 ;
      RECT 179.31 39.34 179.47 43.45 ;
      RECT 179.25 14.84 179.41 16.05 ;
      RECT 179.07 57.79 179.23 62.72 ;
      RECT 177.69 6.24 179.19 6.84 ;
      RECT 178.83 29.97 178.99 32.28 ;
      RECT 178.83 35.23 178.99 36.31 ;
      RECT 178.83 37.11 178.99 38.19 ;
      RECT 178.83 41.14 178.99 43.45 ;
      RECT 178.59 57.79 178.75 62.72 ;
      RECT 178.37 19.63 178.69 20.04 ;
      RECT 178.43 47.88 178.59 51.16 ;
      RECT 177.93 13.8 178.49 13.96 ;
      RECT 177.81 13.32 178.29 13.56 ;
      RECT 178.09 36.21 178.29 36.95 ;
      RECT 178.11 26.38 178.27 27.85 ;
      RECT 178.11 29.32 178.27 34.08 ;
      RECT 178.11 39.34 178.27 46.59 ;
      RECT 178.11 47.59 178.27 51.92 ;
      RECT 178.11 52.64 178.27 56.5 ;
      RECT 177.79 47.88 177.95 51.16 ;
      RECT 177.39 16.47 177.81 17.1 ;
      RECT 177.63 57.79 177.79 62.72 ;
      RECT 177.39 29.97 177.55 32.28 ;
      RECT 177.39 35.23 177.55 36.31 ;
      RECT 177.39 37.11 177.55 38.19 ;
      RECT 177.39 41.14 177.55 43.45 ;
      RECT 177.15 57.79 177.31 62.72 ;
      RECT 176.79 56.99 177.19 57.29 ;
      RECT 176.91 29.97 177.07 34.08 ;
      RECT 176.91 39.34 177.07 43.45 ;
      RECT 176.83 48.24 176.99 50.5 ;
      RECT 176.67 57.79 176.83 67.9 ;
      RECT 174.79 510.54 176.79 510.94 ;
      RECT 176.1 28.33 176.66 28.49 ;
      RECT 176.35 25.51 176.59 26.2 ;
      RECT 176.43 29.97 176.59 32.28 ;
      RECT 176.43 35.23 176.59 36.31 ;
      RECT 176.43 37.11 176.59 38.19 ;
      RECT 176.43 41.14 176.59 43.45 ;
      RECT 175.29 6.24 176.29 6.84 ;
      RECT 175.75 23.54 176.19 23.81 ;
      RECT 175.69 36.21 175.89 36.95 ;
      RECT 175.71 29.32 175.87 34.08 ;
      RECT 175.71 39.34 175.87 46.59 ;
      RECT 175.71 47.59 175.87 51.11 ;
      RECT 175.71 51.34 175.87 53.67 ;
      RECT 175.71 54.16 175.87 56.5 ;
      RECT 175.51 21.85 175.67 22.91 ;
      RECT 175.48 7.58 175.64 8.64 ;
      RECT 175.44 20.65 175.6 21.69 ;
      RECT 174.13 16.8 175.15 17.08 ;
      RECT 174.99 29.97 175.15 32.28 ;
      RECT 174.99 35.23 175.15 36.31 ;
      RECT 174.99 37.11 175.15 38.19 ;
      RECT 174.99 41.14 175.15 43.45 ;
      RECT 174.67 15.32 175.07 15.64 ;
      RECT 174.75 57.79 174.91 67.9 ;
      RECT 174.39 56.99 174.79 57.29 ;
      RECT 174.6 8.04 174.76 8.6 ;
      RECT 174.59 48.24 174.75 50.5 ;
      RECT 174.13 16.12 174.69 16.28 ;
      RECT 174.52 26.68 174.68 28.17 ;
      RECT 174.51 29.97 174.67 34.08 ;
      RECT 174.51 39.34 174.67 43.45 ;
      RECT 174.27 11.52 174.43 13.07 ;
      RECT 174.27 57.79 174.43 62.72 ;
      RECT 174.03 29.97 174.19 32.28 ;
      RECT 174.03 35.23 174.19 36.31 ;
      RECT 174.03 37.11 174.19 38.19 ;
      RECT 174.03 41.14 174.19 43.45 ;
      RECT 173.91 13.11 174.07 13.67 ;
      RECT 173.79 57.79 173.95 62.72 ;
      RECT 172.99 6.24 173.79 6.84 ;
      RECT 173.63 47.88 173.79 51.16 ;
      RECT 173.29 36.21 173.49 36.95 ;
      RECT 173.31 21.45 173.47 24.52 ;
      RECT 173.31 29.32 173.47 34.08 ;
      RECT 173.31 39.34 173.47 46.59 ;
      RECT 173.31 47.59 173.47 51.92 ;
      RECT 173.31 52.64 173.47 56.5 ;
      RECT 172.99 47.88 173.15 51.16 ;
      RECT 172.83 57.79 172.99 62.72 ;
      RECT 172.71 13.11 172.87 13.67 ;
      RECT 172.59 29.97 172.75 32.28 ;
      RECT 172.59 35.23 172.75 36.31 ;
      RECT 172.59 37.11 172.75 38.19 ;
      RECT 172.59 41.14 172.75 43.45 ;
      RECT 172.09 16.12 172.65 16.28 ;
      RECT 171.63 16.8 172.65 17.08 ;
      RECT 172.35 11.52 172.51 13.07 ;
      RECT 172.35 57.79 172.51 62.72 ;
      RECT 171.99 56.99 172.39 57.29 ;
      RECT 172.11 29.97 172.27 34.08 ;
      RECT 172.11 39.34 172.27 43.45 ;
      RECT 172.1 26.68 172.26 28.17 ;
      RECT 172.03 48.24 172.19 50.5 ;
      RECT 172.02 8.04 172.18 8.6 ;
      RECT 171.71 15.32 172.11 15.64 ;
      RECT 171.87 57.79 172.03 67.9 ;
      RECT 169.99 510.54 171.99 510.94 ;
      RECT 171.63 29.97 171.79 32.28 ;
      RECT 171.63 35.23 171.79 36.31 ;
      RECT 171.63 37.11 171.79 38.19 ;
      RECT 171.63 41.14 171.79 43.45 ;
      RECT 170.49 6.24 171.49 6.84 ;
      RECT 171.18 20.65 171.34 21.69 ;
      RECT 171.14 7.58 171.3 8.64 ;
      RECT 171.11 21.85 171.27 22.91 ;
      RECT 170.89 36.21 171.09 36.95 ;
      RECT 170.91 29.32 171.07 34.08 ;
      RECT 170.91 39.34 171.07 46.59 ;
      RECT 170.91 47.59 171.07 51.11 ;
      RECT 170.91 51.34 171.07 53.67 ;
      RECT 170.91 54.16 171.07 56.5 ;
      RECT 170.59 23.54 171.03 23.81 ;
      RECT 170.12 28.33 170.68 28.49 ;
      RECT 170.19 25.51 170.43 26.2 ;
      RECT 170.19 29.97 170.35 32.28 ;
      RECT 170.19 35.23 170.35 36.31 ;
      RECT 170.19 37.11 170.35 38.19 ;
      RECT 170.19 41.14 170.35 43.45 ;
      RECT 169.95 57.79 170.11 67.9 ;
      RECT 169.59 56.99 169.99 57.29 ;
      RECT 169.79 48.24 169.95 50.5 ;
      RECT 169.71 29.97 169.87 34.08 ;
      RECT 169.71 39.34 169.87 43.45 ;
      RECT 169.47 57.79 169.63 62.72 ;
      RECT 168.97 16.47 169.39 17.1 ;
      RECT 169.23 29.97 169.39 32.28 ;
      RECT 169.23 35.23 169.39 36.31 ;
      RECT 169.23 37.11 169.39 38.19 ;
      RECT 169.23 41.14 169.39 43.45 ;
      RECT 168.99 57.79 169.15 62.72 ;
      RECT 167.59 6.24 169.09 6.84 ;
      RECT 168.83 47.88 168.99 51.16 ;
      RECT 168.49 13.32 168.97 13.56 ;
      RECT 168.29 13.8 168.85 13.96 ;
      RECT 168.49 36.21 168.69 36.95 ;
      RECT 168.51 26.38 168.67 27.85 ;
      RECT 168.51 29.32 168.67 34.08 ;
      RECT 168.51 39.34 168.67 46.59 ;
      RECT 168.51 47.59 168.67 51.92 ;
      RECT 168.51 52.64 168.67 56.5 ;
      RECT 168.09 19.63 168.41 20.04 ;
      RECT 168.19 47.88 168.35 51.16 ;
      RECT 168.03 57.79 168.19 62.72 ;
      RECT 167.79 29.97 167.95 32.28 ;
      RECT 167.79 35.23 167.95 36.31 ;
      RECT 167.79 37.11 167.95 38.19 ;
      RECT 167.79 41.14 167.95 43.45 ;
      RECT 167.55 57.79 167.71 62.72 ;
      RECT 167.19 56.99 167.59 57.29 ;
      RECT 167.37 14.84 167.53 16.05 ;
      RECT 167.31 29.97 167.47 34.08 ;
      RECT 167.31 39.34 167.47 43.45 ;
      RECT 167.23 48.24 167.39 50.5 ;
      RECT 167.22 16.21 167.38 18.62 ;
      RECT 167.07 57.79 167.23 67.9 ;
      RECT 165.19 510.54 167.19 510.94 ;
      RECT 165.19 6.24 167.16 6.84 ;
      RECT 166.5 28.33 167.06 28.49 ;
      RECT 166.75 25.51 166.99 26.2 ;
      RECT 166.83 29.97 166.99 32.28 ;
      RECT 166.83 35.23 166.99 36.31 ;
      RECT 166.83 37.11 166.99 38.19 ;
      RECT 166.83 41.14 166.99 43.45 ;
      RECT 166.15 23.54 166.59 23.81 ;
      RECT 166.34 15.33 166.5 15.89 ;
      RECT 166.09 36.21 166.29 36.95 ;
      RECT 166.11 29.32 166.27 34.08 ;
      RECT 166.11 39.34 166.27 46.59 ;
      RECT 166.11 47.59 166.27 51.11 ;
      RECT 166.11 51.34 166.27 53.67 ;
      RECT 166.11 54.16 166.27 56.5 ;
      RECT 164.85 13.4 165.97 13.56 ;
      RECT 165.7 17 165.86 18.12 ;
      RECT 165.05 10 165.77 10.18 ;
      RECT 165.39 29.97 165.55 32.28 ;
      RECT 165.39 35.23 165.55 36.31 ;
      RECT 165.39 37.11 165.55 38.19 ;
      RECT 165.39 41.14 165.55 43.45 ;
      RECT 165.03 10.76 165.35 11.16 ;
      RECT 165.15 57.79 165.31 67.9 ;
      RECT 164.79 56.99 165.19 57.29 ;
      RECT 164.99 48.24 165.15 50.5 ;
      RECT 164.92 26.68 165.08 28.17 ;
      RECT 164.91 29.97 165.07 34.08 ;
      RECT 164.91 39.34 165.07 43.45 ;
      RECT 164.67 57.79 164.83 62.72 ;
      RECT 162.79 6.24 164.79 6.84 ;
      RECT 164.43 29.97 164.59 32.28 ;
      RECT 164.43 35.23 164.59 36.31 ;
      RECT 164.43 37.11 164.59 38.19 ;
      RECT 164.43 41.14 164.59 43.45 ;
      RECT 164.23 12.28 164.55 12.76 ;
      RECT 164.03 8.96 164.54 9.17 ;
      RECT 164.35 21.73 164.51 22.33 ;
      RECT 164.35 22.49 164.51 23.06 ;
      RECT 164.19 57.79 164.35 62.72 ;
      RECT 164.05 15.09 164.33 15.41 ;
      RECT 164.03 47.88 164.19 51.16 ;
      RECT 163.69 36.21 163.89 36.95 ;
      RECT 163.71 21.45 163.87 24.52 ;
      RECT 163.71 29.32 163.87 34.08 ;
      RECT 163.71 39.34 163.87 46.59 ;
      RECT 163.71 47.59 163.87 51.92 ;
      RECT 163.71 52.64 163.87 56.5 ;
      RECT 163.39 47.83 163.55 51.16 ;
      RECT 163.23 57.79 163.39 62.72 ;
      RECT 162.99 29.97 163.15 32.28 ;
      RECT 162.99 35.23 163.15 36.31 ;
      RECT 162.99 37.11 163.15 38.19 ;
      RECT 162.99 41.14 163.15 43.45 ;
      RECT 155.07 15.46 162.91 16.9 ;
      RECT 162.75 57.79 162.91 62.72 ;
      RECT 162.39 56.99 162.79 57.29 ;
      RECT 162.51 29.97 162.67 34.08 ;
      RECT 162.51 39.34 162.67 43.45 ;
      RECT 162.43 48.24 162.59 50.5 ;
      RECT 162.27 57.79 162.43 67.9 ;
      RECT 160.39 510.54 162.39 510.94 ;
      RECT 160.39 6.24 162.37 6.84 ;
      RECT 162.03 29.97 162.19 32.28 ;
      RECT 162.03 35.23 162.19 36.31 ;
      RECT 162.03 37.11 162.19 38.19 ;
      RECT 162.03 41.14 162.19 43.45 ;
      RECT 155.97 21.67 162.01 21.95 ;
      RECT 161.29 36.21 161.49 36.95 ;
      RECT 161.31 29.32 161.47 34.08 ;
      RECT 161.31 39.34 161.47 46.59 ;
      RECT 161.31 47.59 161.47 51.11 ;
      RECT 161.31 51.34 161.47 53.67 ;
      RECT 161.31 54.16 161.47 56.5 ;
      RECT 160.59 29.97 160.75 32.28 ;
      RECT 160.59 35.23 160.75 36.31 ;
      RECT 160.59 37.11 160.75 38.19 ;
      RECT 160.59 41.14 160.75 43.45 ;
      RECT 160.35 57.79 160.51 67.9 ;
      RECT 159.99 56.99 160.39 57.29 ;
      RECT 160.19 48.24 160.35 50.5 ;
      RECT 160.11 29.97 160.27 34.08 ;
      RECT 160.11 39.34 160.27 43.45 ;
      RECT 159.87 57.79 160.03 62.72 ;
      RECT 157.99 6.24 159.97 6.84 ;
      RECT 159.63 29.97 159.79 32.28 ;
      RECT 159.63 35.23 159.79 36.31 ;
      RECT 159.63 37.11 159.79 38.19 ;
      RECT 159.63 41.14 159.79 43.45 ;
      RECT 159.39 57.79 159.55 62.72 ;
      RECT 159.23 47.88 159.39 51.16 ;
      RECT 158.71 9.36 159.27 9.52 ;
      RECT 158.71 11.3 159.27 11.46 ;
      RECT 158.71 14.68 159.27 14.84 ;
      RECT 158.71 19.63 159.27 19.79 ;
      RECT 158.89 36.21 159.09 36.95 ;
      RECT 158.91 29.32 159.07 34.08 ;
      RECT 158.91 39.34 159.07 46.59 ;
      RECT 158.91 47.59 159.07 51.92 ;
      RECT 158.91 52.64 159.07 56.5 ;
      RECT 158.59 47.88 158.75 51.16 ;
      RECT 158.43 57.79 158.59 62.72 ;
      RECT 158.19 29.97 158.35 32.28 ;
      RECT 158.19 35.23 158.35 36.31 ;
      RECT 158.19 37.11 158.35 38.19 ;
      RECT 158.19 41.14 158.35 43.45 ;
      RECT 157.95 57.79 158.11 62.72 ;
      RECT 157.59 56.99 157.99 57.29 ;
      RECT 157.71 29.97 157.87 34.08 ;
      RECT 157.71 39.34 157.87 43.45 ;
      RECT 157.63 48.24 157.79 50.5 ;
      RECT 157.47 57.79 157.63 67.9 ;
      RECT 155.59 510.54 157.59 510.94 ;
      RECT 155.59 6.24 157.57 6.84 ;
      RECT 157.23 29.97 157.39 32.28 ;
      RECT 157.23 35.23 157.39 36.31 ;
      RECT 157.23 37.11 157.39 38.19 ;
      RECT 157.23 41.14 157.39 43.45 ;
      RECT 156.49 36.21 156.69 36.95 ;
      RECT 156.51 29.32 156.67 34.08 ;
      RECT 156.51 39.34 156.67 46.59 ;
      RECT 156.51 47.59 156.67 51.11 ;
      RECT 156.51 51.34 156.67 53.67 ;
      RECT 156.51 54.16 156.67 56.5 ;
      RECT 155.79 29.97 155.95 32.28 ;
      RECT 155.79 35.23 155.95 36.31 ;
      RECT 155.79 37.11 155.95 38.19 ;
      RECT 155.79 41.14 155.95 43.45 ;
      RECT 155.55 57.79 155.71 67.9 ;
      RECT 155.19 56.99 155.59 57.29 ;
      RECT 155.39 48.24 155.55 50.5 ;
      RECT 155.31 29.97 155.47 34.08 ;
      RECT 155.31 39.34 155.47 43.45 ;
      RECT 155.07 57.79 155.23 62.72 ;
      RECT 153.89 6.24 155.19 6.84 ;
      RECT 154.83 29.97 154.99 32.28 ;
      RECT 154.83 35.23 154.99 36.31 ;
      RECT 154.83 37.11 154.99 38.19 ;
      RECT 154.83 41.14 154.99 43.45 ;
      RECT 154.59 57.79 154.75 62.72 ;
      RECT 154.43 47.88 154.59 51.16 ;
      RECT 154.09 36.21 154.29 36.95 ;
      RECT 154.11 29.32 154.27 34.08 ;
      RECT 154.11 39.34 154.27 46.59 ;
      RECT 154.11 47.59 154.27 51.92 ;
      RECT 154.11 52.64 154.27 56.5 ;
      RECT 141.49 7.32 153.69 7.92 ;
      RECT 153.51 63.19 153.67 68.66 ;
      RECT 153.17 57.32 153.33 60.88 ;
      RECT 152.97 32.92 153.13 54.48 ;
      RECT 151.99 510.36 152.79 510.94 ;
      RECT 152.51 51.98 152.67 52.54 ;
      RECT 151.62 44.23 152.02 44.55 ;
      RECT 151.62 44.83 152.02 45.15 ;
      RECT 151.62 45.43 152.02 45.75 ;
      RECT 151.62 46.03 152.02 46.35 ;
      RECT 151.62 46.63 152.02 46.95 ;
      RECT 151.62 47.23 152.02 47.55 ;
      RECT 151.62 47.83 152.02 48.15 ;
      RECT 151.62 48.43 152.02 48.75 ;
      RECT 151.62 49.03 152.02 49.35 ;
      RECT 151.62 49.63 152.02 49.95 ;
      RECT 151.75 22.49 151.91 25.4 ;
      RECT 151.29 6.24 151.89 6.84 ;
      RECT 151.37 22.73 151.59 23.18 ;
      RECT 150.97 54.96 151.13 57.28 ;
      RECT 150.29 6.24 150.89 6.84 ;
      RECT 150.51 43.19 150.67 46.31 ;
      RECT 150.51 48.75 150.67 62.84 ;
      RECT 150.51 63.17 150.67 67.36 ;
      RECT 150.39 30.95 150.55 32.75 ;
      RECT 150.18 69.56 150.4 504.76 ;
      RECT 150.21 29.4 150.37 29.96 ;
      RECT 149.97 52.72 150.25 66.71 ;
      RECT 150.05 27.33 150.21 29.24 ;
      RECT 149.99 22.49 150.15 25.37 ;
      RECT 149.81 29.4 149.97 30.22 ;
      RECT 149.29 35.36 149.97 35.52 ;
      RECT 148.55 22.88 149.83 23.04 ;
      RECT 144.63 69.48 149.77 69.64 ;
      RECT 145.22 70.44 149.77 70.6 ;
      RECT 149.63 70.9 149.77 71.6 ;
      RECT 145.22 71.92 149.77 72.08 ;
      RECT 144.57 72.88 149.77 73.04 ;
      RECT 145.22 73.84 149.77 74 ;
      RECT 149.63 74.32 149.77 75.02 ;
      RECT 145.22 75.32 149.77 75.48 ;
      RECT 144.63 76.28 149.77 76.44 ;
      RECT 145.22 77.24 149.77 77.4 ;
      RECT 149.63 77.7 149.77 78.4 ;
      RECT 145.22 78.72 149.77 78.88 ;
      RECT 144.57 79.68 149.77 79.84 ;
      RECT 145.22 80.64 149.77 80.8 ;
      RECT 149.63 81.12 149.77 81.82 ;
      RECT 145.22 82.12 149.77 82.28 ;
      RECT 144.63 83.08 149.77 83.24 ;
      RECT 145.22 84.04 149.77 84.2 ;
      RECT 149.63 84.5 149.77 85.2 ;
      RECT 145.22 85.52 149.77 85.68 ;
      RECT 144.57 86.48 149.77 86.64 ;
      RECT 145.22 87.44 149.77 87.6 ;
      RECT 149.63 87.92 149.77 88.62 ;
      RECT 145.22 88.92 149.77 89.08 ;
      RECT 144.63 89.88 149.77 90.04 ;
      RECT 145.22 90.84 149.77 91 ;
      RECT 149.63 91.3 149.77 92 ;
      RECT 145.22 92.32 149.77 92.48 ;
      RECT 144.57 93.28 149.77 93.44 ;
      RECT 145.22 94.24 149.77 94.4 ;
      RECT 149.63 94.72 149.77 95.42 ;
      RECT 145.22 95.72 149.77 95.88 ;
      RECT 144.63 96.68 149.77 96.84 ;
      RECT 145.22 97.64 149.77 97.8 ;
      RECT 149.63 98.1 149.77 98.8 ;
      RECT 145.22 99.12 149.77 99.28 ;
      RECT 144.57 100.08 149.77 100.24 ;
      RECT 145.22 101.04 149.77 101.2 ;
      RECT 149.63 101.52 149.77 102.22 ;
      RECT 145.22 102.52 149.77 102.68 ;
      RECT 144.63 103.48 149.77 103.64 ;
      RECT 145.22 104.44 149.77 104.6 ;
      RECT 149.63 104.9 149.77 105.6 ;
      RECT 145.22 105.92 149.77 106.08 ;
      RECT 144.57 106.88 149.77 107.04 ;
      RECT 145.22 107.84 149.77 108 ;
      RECT 149.63 108.32 149.77 109.02 ;
      RECT 145.22 109.32 149.77 109.48 ;
      RECT 144.63 110.28 149.77 110.44 ;
      RECT 145.22 111.24 149.77 111.4 ;
      RECT 149.63 111.7 149.77 112.4 ;
      RECT 145.22 112.72 149.77 112.88 ;
      RECT 144.57 113.68 149.77 113.84 ;
      RECT 145.22 114.64 149.77 114.8 ;
      RECT 149.63 115.12 149.77 115.82 ;
      RECT 145.22 116.12 149.77 116.28 ;
      RECT 144.63 117.08 149.77 117.24 ;
      RECT 145.22 118.04 149.77 118.2 ;
      RECT 149.63 118.5 149.77 119.2 ;
      RECT 145.22 119.52 149.77 119.68 ;
      RECT 144.57 120.48 149.77 120.64 ;
      RECT 145.22 121.44 149.77 121.6 ;
      RECT 149.63 121.92 149.77 122.62 ;
      RECT 145.22 122.92 149.77 123.08 ;
      RECT 144.63 123.88 149.77 124.04 ;
      RECT 145.22 124.84 149.77 125 ;
      RECT 149.63 125.3 149.77 126 ;
      RECT 145.22 126.32 149.77 126.48 ;
      RECT 144.57 127.28 149.77 127.44 ;
      RECT 145.22 128.24 149.77 128.4 ;
      RECT 149.63 128.72 149.77 129.42 ;
      RECT 145.22 129.72 149.77 129.88 ;
      RECT 144.63 130.68 149.77 130.84 ;
      RECT 145.22 131.64 149.77 131.8 ;
      RECT 149.63 132.1 149.77 132.8 ;
      RECT 145.22 133.12 149.77 133.28 ;
      RECT 144.57 134.08 149.77 134.24 ;
      RECT 145.22 135.04 149.77 135.2 ;
      RECT 149.63 135.52 149.77 136.22 ;
      RECT 145.22 136.52 149.77 136.68 ;
      RECT 144.63 137.48 149.77 137.64 ;
      RECT 145.22 138.44 149.77 138.6 ;
      RECT 149.63 138.9 149.77 139.6 ;
      RECT 145.22 139.92 149.77 140.08 ;
      RECT 144.57 140.88 149.77 141.04 ;
      RECT 145.22 141.84 149.77 142 ;
      RECT 149.63 142.32 149.77 143.02 ;
      RECT 145.22 143.32 149.77 143.48 ;
      RECT 144.63 144.28 149.77 144.44 ;
      RECT 145.22 145.24 149.77 145.4 ;
      RECT 149.63 145.7 149.77 146.4 ;
      RECT 145.22 146.72 149.77 146.88 ;
      RECT 144.57 147.68 149.77 147.84 ;
      RECT 145.22 148.64 149.77 148.8 ;
      RECT 149.63 149.12 149.77 149.82 ;
      RECT 145.22 150.12 149.77 150.28 ;
      RECT 144.63 151.08 149.77 151.24 ;
      RECT 145.22 152.04 149.77 152.2 ;
      RECT 149.63 152.5 149.77 153.2 ;
      RECT 145.22 153.52 149.77 153.68 ;
      RECT 149.55 52.83 149.71 61.96 ;
      RECT 149.55 62.12 149.71 63.79 ;
      RECT 149.55 63.97 149.71 67.36 ;
      RECT 149.21 27.73 149.37 29.28 ;
      RECT 148.01 510.36 149.33 510.94 ;
      RECT 149.01 52.72 149.29 66.71 ;
      RECT 147.89 508.32 148.97 508.48 ;
      RECT 148.01 6.24 148.87 6.84 ;
      RECT 148.53 29.89 148.83 30.45 ;
      RECT 148.59 47.62 148.75 62.84 ;
      RECT 148.59 63.17 148.75 67.36 ;
      RECT 148.41 27.81 148.57 29.3 ;
      RECT 148.35 506.86 148.51 507.94 ;
      RECT 148.23 22.5 148.39 25.37 ;
      RECT 148.05 52.72 148.33 66.71 ;
      RECT 147.37 35.36 148.05 35.52 ;
      RECT 147.79 29.78 147.95 30.47 ;
      RECT 147.63 52.83 147.79 61.96 ;
      RECT 147.63 62.12 147.79 63.79 ;
      RECT 147.63 63.97 147.79 67.36 ;
      RECT 146.85 29.53 147.45 29.73 ;
      RECT 146.09 6.24 147.41 6.84 ;
      RECT 147.09 52.72 147.37 66.71 ;
      RECT 146.15 508.32 147.23 508.48 ;
      RECT 146.33 29.95 147.05 30.11 ;
      RECT 146.67 43.19 146.83 46.31 ;
      RECT 146.67 48.75 146.83 62.84 ;
      RECT 146.67 63.17 146.83 67.36 ;
      RECT 146.59 506.92 146.79 507.94 ;
      RECT 146.59 508.86 146.79 509.88 ;
      RECT 146.49 30.63 146.65 32.41 ;
      RECT 146.47 22.5 146.63 25.37 ;
      RECT 146.13 52.72 146.41 66.71 ;
      RECT 146.03 22.38 146.27 23.12 ;
      RECT 146.08 14.87 146.24 17.13 ;
      RECT 145.45 35.36 146.13 35.52 ;
      RECT 145.36 15.97 145.92 16.13 ;
      RECT 145.71 52.83 145.87 61.96 ;
      RECT 145.71 62.12 145.87 63.79 ;
      RECT 145.71 63.97 145.87 67.36 ;
      RECT 145.49 30.63 145.65 32.53 ;
      RECT 145.01 6.24 145.61 6.84 ;
      RECT 144.41 508.32 145.49 508.48 ;
      RECT 144.17 510.36 145.49 510.94 ;
      RECT 145.17 52.72 145.45 66.71 ;
      RECT 144.85 506.92 145.05 507.94 ;
      RECT 144.85 508.86 145.05 509.88 ;
      RECT 144.75 47.62 144.91 62.84 ;
      RECT 144.75 63.17 144.91 67.36 ;
      RECT 144.67 29.6 144.85 30.67 ;
      RECT 143.94 505.84 144.66 506 ;
      RECT 144.49 16.08 144.65 16.64 ;
      RECT 144.21 52.72 144.49 66.71 ;
      RECT 144.17 15.66 144.33 17.4 ;
      RECT 143.53 35.36 144.21 35.52 ;
      RECT 143.9 30.63 144.06 32.25 ;
      RECT 131.27 69.48 143.97 69.64 ;
      RECT 131.27 72.88 143.97 73.04 ;
      RECT 131.27 76.28 143.97 76.44 ;
      RECT 131.27 79.68 143.97 79.84 ;
      RECT 131.27 83.08 143.97 83.24 ;
      RECT 131.27 86.48 143.97 86.64 ;
      RECT 131.27 89.88 143.97 90.04 ;
      RECT 131.27 93.28 143.97 93.44 ;
      RECT 131.27 96.68 143.97 96.84 ;
      RECT 131.27 100.08 143.97 100.24 ;
      RECT 131.27 103.48 143.97 103.64 ;
      RECT 131.27 106.88 143.97 107.04 ;
      RECT 131.27 110.28 143.97 110.44 ;
      RECT 131.27 113.68 143.97 113.84 ;
      RECT 131.27 117.08 143.97 117.24 ;
      RECT 131.27 120.48 143.97 120.64 ;
      RECT 131.27 123.88 143.97 124.04 ;
      RECT 131.27 127.28 143.97 127.44 ;
      RECT 131.27 130.68 143.97 130.84 ;
      RECT 131.27 134.08 143.97 134.24 ;
      RECT 131.27 137.48 143.97 137.64 ;
      RECT 131.27 140.88 143.97 141.04 ;
      RECT 131.27 144.28 143.97 144.44 ;
      RECT 131.27 147.68 143.97 147.84 ;
      RECT 131.27 151.08 143.97 151.24 ;
      RECT 131.27 154.48 143.97 154.64 ;
      RECT 131.27 157.88 143.97 158.04 ;
      RECT 131.27 161.28 143.97 161.44 ;
      RECT 131.27 164.68 143.97 164.84 ;
      RECT 131.27 168.08 143.97 168.24 ;
      RECT 131.27 171.48 143.97 171.64 ;
      RECT 131.27 174.88 143.97 175.04 ;
      RECT 131.27 178.28 143.97 178.44 ;
      RECT 131.27 181.68 143.97 181.84 ;
      RECT 131.27 185.08 143.97 185.24 ;
      RECT 131.27 188.48 143.97 188.64 ;
      RECT 131.27 191.88 143.97 192.04 ;
      RECT 131.27 195.28 143.97 195.44 ;
      RECT 131.27 198.68 143.97 198.84 ;
      RECT 131.27 202.08 143.97 202.24 ;
      RECT 131.27 205.48 143.97 205.64 ;
      RECT 131.27 208.88 143.97 209.04 ;
      RECT 131.27 212.28 143.97 212.44 ;
      RECT 131.27 215.68 143.97 215.84 ;
      RECT 131.27 219.08 143.97 219.24 ;
      RECT 131.27 222.48 143.97 222.64 ;
      RECT 131.27 225.88 143.97 226.04 ;
      RECT 131.27 229.28 143.97 229.44 ;
      RECT 131.27 232.68 143.97 232.84 ;
      RECT 131.27 236.08 143.97 236.24 ;
      RECT 131.27 239.48 143.97 239.64 ;
      RECT 131.27 242.88 143.97 243.04 ;
      RECT 131.27 246.28 143.97 246.44 ;
      RECT 131.27 249.68 143.97 249.84 ;
      RECT 131.27 253.08 143.97 253.24 ;
      RECT 131.27 256.48 143.97 256.64 ;
      RECT 131.27 259.88 143.97 260.04 ;
      RECT 131.27 263.28 143.97 263.44 ;
      RECT 131.27 266.68 143.97 266.84 ;
      RECT 131.27 270.08 143.97 270.24 ;
      RECT 131.27 273.48 143.97 273.64 ;
      RECT 131.27 276.88 143.97 277.04 ;
      RECT 131.27 280.28 143.97 280.44 ;
      RECT 131.27 283.68 143.97 283.84 ;
      RECT 131.27 287.08 143.97 287.24 ;
      RECT 131.27 290.48 143.97 290.64 ;
      RECT 131.27 293.88 143.97 294.04 ;
      RECT 131.27 297.28 143.97 297.44 ;
      RECT 131.27 300.68 143.97 300.84 ;
      RECT 131.27 304.08 143.97 304.24 ;
      RECT 131.27 307.48 143.97 307.64 ;
      RECT 131.27 310.88 143.97 311.04 ;
      RECT 131.27 314.28 143.97 314.44 ;
      RECT 131.27 317.68 143.97 317.84 ;
      RECT 131.27 321.08 143.97 321.24 ;
      RECT 131.27 324.48 143.97 324.64 ;
      RECT 131.27 327.88 143.97 328.04 ;
      RECT 131.27 331.28 143.97 331.44 ;
      RECT 131.27 334.68 143.97 334.84 ;
      RECT 131.27 338.08 143.97 338.24 ;
      RECT 131.27 341.48 143.97 341.64 ;
      RECT 131.27 344.88 143.97 345.04 ;
      RECT 131.27 348.28 143.97 348.44 ;
      RECT 131.27 351.68 143.97 351.84 ;
      RECT 131.27 355.08 143.97 355.24 ;
      RECT 131.27 358.48 143.97 358.64 ;
      RECT 131.27 361.88 143.97 362.04 ;
      RECT 131.27 365.28 143.97 365.44 ;
      RECT 131.27 368.68 143.97 368.84 ;
      RECT 131.27 372.08 143.97 372.24 ;
      RECT 131.27 375.48 143.97 375.64 ;
      RECT 131.27 378.88 143.97 379.04 ;
      RECT 131.27 382.28 143.97 382.44 ;
      RECT 131.27 385.68 143.97 385.84 ;
      RECT 131.27 389.08 143.97 389.24 ;
      RECT 131.27 392.48 143.97 392.64 ;
      RECT 131.27 395.88 143.97 396.04 ;
      RECT 131.27 399.28 143.97 399.44 ;
      RECT 131.27 402.68 143.97 402.84 ;
      RECT 131.27 406.08 143.97 406.24 ;
      RECT 131.27 409.48 143.97 409.64 ;
      RECT 131.27 412.88 143.97 413.04 ;
      RECT 131.27 416.28 143.97 416.44 ;
      RECT 131.27 419.68 143.97 419.84 ;
      RECT 131.27 423.08 143.97 423.24 ;
      RECT 131.27 426.48 143.97 426.64 ;
      RECT 131.27 429.88 143.97 430.04 ;
      RECT 131.27 433.28 143.97 433.44 ;
      RECT 131.27 436.68 143.97 436.84 ;
      RECT 131.27 440.08 143.97 440.24 ;
      RECT 131.27 443.48 143.97 443.64 ;
      RECT 131.27 446.88 143.97 447.04 ;
      RECT 131.27 450.28 143.97 450.44 ;
      RECT 131.27 453.68 143.97 453.84 ;
      RECT 131.27 457.08 143.97 457.24 ;
      RECT 131.27 460.48 143.97 460.64 ;
      RECT 131.27 463.88 143.97 464.04 ;
      RECT 131.27 467.28 143.97 467.44 ;
      RECT 131.27 470.68 143.97 470.84 ;
      RECT 131.27 474.08 143.97 474.24 ;
      RECT 131.27 477.48 143.97 477.64 ;
      RECT 131.27 480.88 143.97 481.04 ;
      RECT 131.27 484.28 143.97 484.44 ;
      RECT 131.27 487.68 143.97 487.84 ;
      RECT 131.27 491.08 143.97 491.24 ;
      RECT 131.27 494.48 143.97 494.64 ;
      RECT 131.27 497.88 143.97 498.04 ;
      RECT 131.27 501.28 143.97 501.44 ;
      RECT 143.79 52.83 143.95 61.96 ;
      RECT 143.79 62.12 143.95 63.79 ;
      RECT 143.79 63.97 143.95 67.36 ;
      RECT 142.67 508.32 143.75 508.48 ;
      RECT 143.25 52.72 143.53 66.71 ;
      RECT 143.26 30.13 143.42 30.74 ;
      RECT 135.81 70.44 143.38 70.6 ;
      RECT 135.8 71.92 143.38 72.08 ;
      RECT 135.8 73.84 143.38 74 ;
      RECT 135.81 75.32 143.38 75.48 ;
      RECT 135.81 77.24 143.38 77.4 ;
      RECT 135.8 78.72 143.38 78.88 ;
      RECT 135.8 80.64 143.38 80.8 ;
      RECT 135.81 82.12 143.38 82.28 ;
      RECT 135.81 84.04 143.38 84.2 ;
      RECT 135.8 85.52 143.38 85.68 ;
      RECT 135.8 87.44 143.38 87.6 ;
      RECT 135.81 88.92 143.38 89.08 ;
      RECT 135.81 90.84 143.38 91 ;
      RECT 135.8 92.32 143.38 92.48 ;
      RECT 135.8 94.24 143.38 94.4 ;
      RECT 135.81 95.72 143.38 95.88 ;
      RECT 135.81 97.64 143.38 97.8 ;
      RECT 135.8 99.12 143.38 99.28 ;
      RECT 135.8 101.04 143.38 101.2 ;
      RECT 135.81 102.52 143.38 102.68 ;
      RECT 135.81 104.44 143.38 104.6 ;
      RECT 135.8 105.92 143.38 106.08 ;
      RECT 135.8 107.84 143.38 108 ;
      RECT 135.81 109.32 143.38 109.48 ;
      RECT 135.81 111.24 143.38 111.4 ;
      RECT 135.8 112.72 143.38 112.88 ;
      RECT 135.8 114.64 143.38 114.8 ;
      RECT 135.81 116.12 143.38 116.28 ;
      RECT 135.81 118.04 143.38 118.2 ;
      RECT 135.8 119.52 143.38 119.68 ;
      RECT 135.8 121.44 143.38 121.6 ;
      RECT 135.81 122.92 143.38 123.08 ;
      RECT 135.81 124.84 143.38 125 ;
      RECT 135.8 126.32 143.38 126.48 ;
      RECT 135.8 128.24 143.38 128.4 ;
      RECT 135.81 129.72 143.38 129.88 ;
      RECT 135.81 131.64 143.38 131.8 ;
      RECT 135.8 133.12 143.38 133.28 ;
      RECT 135.8 135.04 143.38 135.2 ;
      RECT 135.81 136.52 143.38 136.68 ;
      RECT 135.81 138.44 143.38 138.6 ;
      RECT 135.8 139.92 143.38 140.08 ;
      RECT 135.8 141.84 143.38 142 ;
      RECT 135.81 143.32 143.38 143.48 ;
      RECT 135.81 145.24 143.38 145.4 ;
      RECT 135.8 146.72 143.38 146.88 ;
      RECT 135.8 148.64 143.38 148.8 ;
      RECT 135.81 150.12 143.38 150.28 ;
      RECT 135.81 152.04 143.38 152.2 ;
      RECT 135.8 153.52 143.38 153.68 ;
      RECT 135.8 155.44 143.38 155.6 ;
      RECT 135.81 156.92 143.38 157.08 ;
      RECT 135.81 158.84 143.38 159 ;
      RECT 135.8 160.32 143.38 160.48 ;
      RECT 135.8 162.24 143.38 162.4 ;
      RECT 135.81 163.72 143.38 163.88 ;
      RECT 135.81 165.64 143.38 165.8 ;
      RECT 135.8 167.12 143.38 167.28 ;
      RECT 135.8 169.04 143.38 169.2 ;
      RECT 135.81 170.52 143.38 170.68 ;
      RECT 135.81 172.44 143.38 172.6 ;
      RECT 135.8 173.92 143.38 174.08 ;
      RECT 135.8 175.84 143.38 176 ;
      RECT 135.81 177.32 143.38 177.48 ;
      RECT 135.81 179.24 143.38 179.4 ;
      RECT 135.8 180.72 143.38 180.88 ;
      RECT 135.8 182.64 143.38 182.8 ;
      RECT 135.81 184.12 143.38 184.28 ;
      RECT 135.81 186.04 143.38 186.2 ;
      RECT 135.8 187.52 143.38 187.68 ;
      RECT 135.8 189.44 143.38 189.6 ;
      RECT 135.81 190.92 143.38 191.08 ;
      RECT 135.81 192.84 143.38 193 ;
      RECT 135.8 194.32 143.38 194.48 ;
      RECT 135.8 196.24 143.38 196.4 ;
      RECT 135.81 197.72 143.38 197.88 ;
      RECT 135.81 199.64 143.38 199.8 ;
      RECT 135.8 201.12 143.38 201.28 ;
      RECT 135.8 203.04 143.38 203.2 ;
      RECT 135.81 204.52 143.38 204.68 ;
      RECT 135.81 206.44 143.38 206.6 ;
      RECT 135.8 207.92 143.38 208.08 ;
      RECT 135.8 209.84 143.38 210 ;
      RECT 135.81 211.32 143.38 211.48 ;
      RECT 135.81 213.24 143.38 213.4 ;
      RECT 135.8 214.72 143.38 214.88 ;
      RECT 135.8 216.64 143.38 216.8 ;
      RECT 135.81 218.12 143.38 218.28 ;
      RECT 135.81 220.04 143.38 220.2 ;
      RECT 135.8 221.52 143.38 221.68 ;
      RECT 135.8 223.44 143.38 223.6 ;
      RECT 135.81 224.92 143.38 225.08 ;
      RECT 135.81 226.84 143.38 227 ;
      RECT 135.8 228.32 143.38 228.48 ;
      RECT 135.8 230.24 143.38 230.4 ;
      RECT 135.81 231.72 143.38 231.88 ;
      RECT 135.81 233.64 143.38 233.8 ;
      RECT 135.8 235.12 143.38 235.28 ;
      RECT 135.8 237.04 143.38 237.2 ;
      RECT 135.81 238.52 143.38 238.68 ;
      RECT 135.81 240.44 143.38 240.6 ;
      RECT 135.8 241.92 143.38 242.08 ;
      RECT 135.8 243.84 143.38 244 ;
      RECT 135.81 245.32 143.38 245.48 ;
      RECT 135.81 247.24 143.38 247.4 ;
      RECT 135.8 248.72 143.38 248.88 ;
      RECT 135.8 250.64 143.38 250.8 ;
      RECT 135.81 252.12 143.38 252.28 ;
      RECT 135.81 254.04 143.38 254.2 ;
      RECT 135.8 255.52 143.38 255.68 ;
      RECT 135.8 257.44 143.38 257.6 ;
      RECT 135.81 258.92 143.38 259.08 ;
      RECT 135.81 260.84 143.38 261 ;
      RECT 135.8 262.32 143.38 262.48 ;
      RECT 135.8 264.24 143.38 264.4 ;
      RECT 135.81 265.72 143.38 265.88 ;
      RECT 135.81 267.64 143.38 267.8 ;
      RECT 135.8 269.12 143.38 269.28 ;
      RECT 135.8 271.04 143.38 271.2 ;
      RECT 135.81 272.52 143.38 272.68 ;
      RECT 135.81 274.44 143.38 274.6 ;
      RECT 135.8 275.92 143.38 276.08 ;
      RECT 135.8 277.84 143.38 278 ;
      RECT 135.81 279.32 143.38 279.48 ;
      RECT 135.81 281.24 143.38 281.4 ;
      RECT 135.8 282.72 143.38 282.88 ;
      RECT 135.8 284.64 143.38 284.8 ;
      RECT 135.81 286.12 143.38 286.28 ;
      RECT 135.81 288.04 143.38 288.2 ;
      RECT 135.8 289.52 143.38 289.68 ;
      RECT 135.8 291.44 143.38 291.6 ;
      RECT 135.81 292.92 143.38 293.08 ;
      RECT 135.81 294.84 143.38 295 ;
      RECT 135.8 296.32 143.38 296.48 ;
      RECT 135.8 298.24 143.38 298.4 ;
      RECT 135.81 299.72 143.38 299.88 ;
      RECT 135.81 301.64 143.38 301.8 ;
      RECT 135.8 303.12 143.38 303.28 ;
      RECT 135.8 305.04 143.38 305.2 ;
      RECT 135.81 306.52 143.38 306.68 ;
      RECT 135.81 308.44 143.38 308.6 ;
      RECT 135.8 309.92 143.38 310.08 ;
      RECT 135.8 311.84 143.38 312 ;
      RECT 135.81 313.32 143.38 313.48 ;
      RECT 135.81 315.24 143.38 315.4 ;
      RECT 135.8 316.72 143.38 316.88 ;
      RECT 135.8 318.64 143.38 318.8 ;
      RECT 135.81 320.12 143.38 320.28 ;
      RECT 135.81 322.04 143.38 322.2 ;
      RECT 135.8 323.52 143.38 323.68 ;
      RECT 135.8 325.44 143.38 325.6 ;
      RECT 135.81 326.92 143.38 327.08 ;
      RECT 135.81 328.84 143.38 329 ;
      RECT 135.8 330.32 143.38 330.48 ;
      RECT 135.8 332.24 143.38 332.4 ;
      RECT 135.81 333.72 143.38 333.88 ;
      RECT 135.81 335.64 143.38 335.8 ;
      RECT 135.8 337.12 143.38 337.28 ;
      RECT 135.8 339.04 143.38 339.2 ;
      RECT 135.81 340.52 143.38 340.68 ;
      RECT 135.81 342.44 143.38 342.6 ;
      RECT 135.8 343.92 143.38 344.08 ;
      RECT 135.8 345.84 143.38 346 ;
      RECT 135.81 347.32 143.38 347.48 ;
      RECT 135.81 349.24 143.38 349.4 ;
      RECT 135.8 350.72 143.38 350.88 ;
      RECT 135.8 352.64 143.38 352.8 ;
      RECT 135.81 354.12 143.38 354.28 ;
      RECT 135.81 356.04 143.38 356.2 ;
      RECT 135.8 357.52 143.38 357.68 ;
      RECT 135.8 359.44 143.38 359.6 ;
      RECT 135.81 360.92 143.38 361.08 ;
      RECT 135.81 362.84 143.38 363 ;
      RECT 135.8 364.32 143.38 364.48 ;
      RECT 135.8 366.24 143.38 366.4 ;
      RECT 135.81 367.72 143.38 367.88 ;
      RECT 135.81 369.64 143.38 369.8 ;
      RECT 135.8 371.12 143.38 371.28 ;
      RECT 135.8 373.04 143.38 373.2 ;
      RECT 135.81 374.52 143.38 374.68 ;
      RECT 135.81 376.44 143.38 376.6 ;
      RECT 135.8 377.92 143.38 378.08 ;
      RECT 135.8 379.84 143.38 380 ;
      RECT 135.81 381.32 143.38 381.48 ;
      RECT 135.81 383.24 143.38 383.4 ;
      RECT 135.8 384.72 143.38 384.88 ;
      RECT 135.8 386.64 143.38 386.8 ;
      RECT 135.81 388.12 143.38 388.28 ;
      RECT 135.81 390.04 143.38 390.2 ;
      RECT 135.8 391.52 143.38 391.68 ;
      RECT 135.8 393.44 143.38 393.6 ;
      RECT 135.81 394.92 143.38 395.08 ;
      RECT 135.81 396.84 143.38 397 ;
      RECT 135.8 398.32 143.38 398.48 ;
      RECT 135.8 400.24 143.38 400.4 ;
      RECT 135.81 401.72 143.38 401.88 ;
      RECT 135.81 403.64 143.38 403.8 ;
      RECT 135.8 405.12 143.38 405.28 ;
      RECT 135.8 407.04 143.38 407.2 ;
      RECT 135.81 408.52 143.38 408.68 ;
      RECT 135.81 410.44 143.38 410.6 ;
      RECT 135.8 411.92 143.38 412.08 ;
      RECT 135.8 413.84 143.38 414 ;
      RECT 135.81 415.32 143.38 415.48 ;
      RECT 135.81 417.24 143.38 417.4 ;
      RECT 135.8 418.72 143.38 418.88 ;
      RECT 135.8 420.64 143.38 420.8 ;
      RECT 135.81 422.12 143.38 422.28 ;
      RECT 135.81 424.04 143.38 424.2 ;
      RECT 135.8 425.52 143.38 425.68 ;
      RECT 135.8 427.44 143.38 427.6 ;
      RECT 135.81 428.92 143.38 429.08 ;
      RECT 135.81 430.84 143.38 431 ;
      RECT 135.8 432.32 143.38 432.48 ;
      RECT 135.8 434.24 143.38 434.4 ;
      RECT 135.81 435.72 143.38 435.88 ;
      RECT 135.81 437.64 143.38 437.8 ;
      RECT 135.8 439.12 143.38 439.28 ;
      RECT 135.8 441.04 143.38 441.2 ;
      RECT 135.81 442.52 143.38 442.68 ;
      RECT 135.81 444.44 143.38 444.6 ;
      RECT 135.8 445.92 143.38 446.08 ;
      RECT 135.8 447.84 143.38 448 ;
      RECT 135.81 449.32 143.38 449.48 ;
      RECT 135.81 451.24 143.38 451.4 ;
      RECT 135.8 452.72 143.38 452.88 ;
      RECT 135.8 454.64 143.38 454.8 ;
      RECT 135.81 456.12 143.38 456.28 ;
      RECT 135.81 458.04 143.38 458.2 ;
      RECT 135.8 459.52 143.38 459.68 ;
      RECT 135.8 461.44 143.38 461.6 ;
      RECT 135.81 462.92 143.38 463.08 ;
      RECT 135.81 464.84 143.38 465 ;
      RECT 135.8 466.32 143.38 466.48 ;
      RECT 135.8 468.24 143.38 468.4 ;
      RECT 135.81 469.72 143.38 469.88 ;
      RECT 135.81 471.64 143.38 471.8 ;
      RECT 135.8 473.12 143.38 473.28 ;
      RECT 135.8 475.04 143.38 475.2 ;
      RECT 135.81 476.52 143.38 476.68 ;
      RECT 135.81 478.44 143.38 478.6 ;
      RECT 135.8 479.92 143.38 480.08 ;
      RECT 135.8 481.84 143.38 482 ;
      RECT 135.81 483.32 143.38 483.48 ;
      RECT 135.81 485.24 143.38 485.4 ;
      RECT 135.8 486.72 143.38 486.88 ;
      RECT 135.8 488.64 143.38 488.8 ;
      RECT 135.81 490.12 143.38 490.28 ;
      RECT 135.81 492.04 143.38 492.2 ;
      RECT 135.8 493.52 143.38 493.68 ;
      RECT 135.8 495.44 143.38 495.6 ;
      RECT 135.81 496.92 143.38 497.08 ;
      RECT 135.81 498.84 143.38 499 ;
      RECT 135.8 500.32 143.38 500.48 ;
      RECT 135.8 502.24 143.38 502.4 ;
      RECT 135.81 503.72 143.38 503.88 ;
      RECT 143.11 506.92 143.31 508 ;
      RECT 143.11 508.8 143.31 509.88 ;
      RECT 142.83 43.19 142.99 46.31 ;
      RECT 142.83 48.75 142.99 62.84 ;
      RECT 142.83 63.17 142.99 67.36 ;
      RECT 142.34 29.66 142.78 29.94 ;
      RECT 142.29 52.72 142.57 66.71 ;
      RECT 141.75 30.1 142.36 30.29 ;
      RECT 141.61 35.36 142.29 35.52 ;
      RECT 141.62 6.24 142.22 6.84 ;
      RECT 141.87 52.83 142.03 61.96 ;
      RECT 141.87 62.12 142.03 63.79 ;
      RECT 141.87 63.97 142.03 67.36 ;
      RECT 140.93 508.32 142.01 508.48 ;
      RECT 138.41 510.54 141.65 510.94 ;
      RECT 141.33 52.72 141.61 66.71 ;
      RECT 141.37 506.92 141.57 508 ;
      RECT 141.37 508.8 141.57 509.88 ;
      RECT 140.91 47.62 141.07 62.84 ;
      RECT 140.91 63.17 141.07 67.36 ;
      RECT 138.83 6.24 140.83 6.84 ;
      RECT 140.51 35.22 140.67 36.23 ;
      RECT 139.19 508.32 140.27 508.48 ;
      RECT 139.71 23.97 139.92 24.48 ;
      RECT 139.7 57.58 139.92 58.08 ;
      RECT 139.73 12.63 139.89 17.44 ;
      RECT 139.73 31.09 139.89 36.97 ;
      RECT 139.73 40.73 139.89 41.55 ;
      RECT 139.73 45.65 139.89 51.3 ;
      RECT 139.63 506.92 139.83 508 ;
      RECT 139.63 508.8 139.83 509.88 ;
      RECT 139.25 9.61 139.41 14.44 ;
      RECT 138.94 37.58 139.23 38.41 ;
      RECT 138.99 30.54 139.15 32.2 ;
      RECT 138.99 50.09 139.15 51.7 ;
      RECT 138.91 38.57 139.07 40.5 ;
      RECT 138.5 37.58 138.78 38.41 ;
      RECT 138.51 17.46 138.67 20.88 ;
      RECT 138.51 61.17 138.67 64.59 ;
      RECT 137.45 508.32 138.53 508.48 ;
      RECT 137.77 23.99 138.45 24.21 ;
      RECT 137.77 57.84 138.45 58.06 ;
      RECT 137.96 7.04 138.28 7.36 ;
      RECT 137.89 506.92 138.09 508 ;
      RECT 137.89 508.8 138.09 509.78 ;
      RECT 137.55 17.46 137.71 20.88 ;
      RECT 137.55 61.17 137.71 64.59 ;
      RECT 137.43 37.58 137.6 38.41 ;
      RECT 135.43 6.24 137.39 6.84 ;
      RECT 137.15 38.57 137.31 40.5 ;
      RECT 136.99 37.58 137.18 38.41 ;
      RECT 136.81 9.61 136.97 14.44 ;
      RECT 136.33 12.63 136.49 17.44 ;
      RECT 136.33 17.6 136.49 20.88 ;
      RECT 136.33 32.85 136.49 36.97 ;
      RECT 136.33 40.73 136.49 41.55 ;
      RECT 136.33 60.41 136.49 64 ;
      RECT 135.85 9.61 136.01 14.44 ;
      RECT 135.64 37.58 135.83 38.41 ;
      RECT 135.51 38.57 135.67 40.5 ;
      RECT 135.22 37.58 135.39 38.41 ;
      RECT 135.11 17.46 135.27 20.88 ;
      RECT 135.11 61.17 135.27 64.59 ;
      RECT 134.37 23.99 135.05 24.21 ;
      RECT 134.37 57.84 135.05 58.06 ;
      RECT 134.54 7.04 134.86 7.36 ;
      RECT 131.61 510.54 134.41 510.94 ;
      RECT 134.04 37.58 134.32 38.41 ;
      RECT 134.15 17.46 134.31 20.88 ;
      RECT 134.15 61.17 134.31 64.59 ;
      RECT 132.03 6.24 133.99 6.84 ;
      RECT 133.75 38.57 133.91 40.5 ;
      RECT 133.59 37.58 133.88 38.41 ;
      RECT 133.67 30.54 133.83 32.2 ;
      RECT 133.67 50.09 133.83 51.7 ;
      RECT 133.41 9.61 133.57 14.44 ;
      RECT 132.9 23.97 133.12 24.48 ;
      RECT 132.9 57.58 133.12 58.08 ;
      RECT 132.93 12.63 133.09 17.44 ;
      RECT 132.93 31.09 133.09 36.97 ;
      RECT 132.93 40.73 133.09 41.55 ;
      RECT 132.93 45.65 133.09 51.3 ;
      RECT 132.45 9.61 132.61 14.44 ;
      RECT 132.14 37.58 132.43 38.41 ;
      RECT 132.19 30.54 132.35 32.2 ;
      RECT 132.19 50.09 132.35 51.7 ;
      RECT 132.11 38.57 132.27 40.5 ;
      RECT 131.7 37.58 131.98 38.41 ;
      RECT 131.71 17.46 131.87 20.88 ;
      RECT 131.71 61.17 131.87 64.59 ;
      RECT 130.97 23.99 131.65 24.21 ;
      RECT 130.97 57.84 131.65 58.06 ;
      RECT 131.16 7.04 131.48 7.36 ;
      RECT 130.75 17.46 130.91 20.88 ;
      RECT 130.75 61.17 130.91 64.59 ;
      RECT 130.63 37.58 130.8 38.41 ;
      RECT 128.63 6.24 130.59 6.84 ;
      RECT 130.35 38.57 130.51 40.5 ;
      RECT 130.19 37.58 130.38 38.41 ;
      RECT 130.01 9.61 130.17 14.44 ;
      RECT 123.49 69.48 129.98 69.64 ;
      RECT 123.47 72.88 129.98 73.04 ;
      RECT 123.49 76.28 129.98 76.44 ;
      RECT 123.47 79.68 129.98 79.84 ;
      RECT 123.49 83.08 129.98 83.24 ;
      RECT 123.47 86.48 129.98 86.64 ;
      RECT 123.49 89.88 129.98 90.04 ;
      RECT 123.47 93.28 129.98 93.44 ;
      RECT 123.49 96.68 129.98 96.84 ;
      RECT 123.47 100.08 129.98 100.24 ;
      RECT 123.49 103.48 129.98 103.64 ;
      RECT 123.47 106.88 129.98 107.04 ;
      RECT 123.49 110.28 129.98 110.44 ;
      RECT 123.47 113.68 129.98 113.84 ;
      RECT 123.49 117.08 129.98 117.24 ;
      RECT 123.47 120.48 129.98 120.64 ;
      RECT 123.49 123.88 129.98 124.04 ;
      RECT 123.47 127.28 129.98 127.44 ;
      RECT 123.49 130.68 129.98 130.84 ;
      RECT 123.47 134.08 129.98 134.24 ;
      RECT 123.49 137.48 129.98 137.64 ;
      RECT 123.47 140.88 129.98 141.04 ;
      RECT 123.49 144.28 129.98 144.44 ;
      RECT 123.47 147.68 129.98 147.84 ;
      RECT 123.49 151.08 129.98 151.24 ;
      RECT 123.47 154.48 129.98 154.64 ;
      RECT 123.49 157.88 129.98 158.04 ;
      RECT 123.47 161.28 129.98 161.44 ;
      RECT 123.49 164.68 129.98 164.84 ;
      RECT 123.47 168.08 129.98 168.24 ;
      RECT 123.49 171.48 129.98 171.64 ;
      RECT 123.47 174.88 129.98 175.04 ;
      RECT 123.49 178.28 129.98 178.44 ;
      RECT 123.47 181.68 129.98 181.84 ;
      RECT 123.49 185.08 129.98 185.24 ;
      RECT 123.47 188.48 129.98 188.64 ;
      RECT 123.49 191.88 129.98 192.04 ;
      RECT 123.47 195.28 129.98 195.44 ;
      RECT 123.49 198.68 129.98 198.84 ;
      RECT 123.47 202.08 129.98 202.24 ;
      RECT 123.49 205.48 129.98 205.64 ;
      RECT 123.47 208.88 129.98 209.04 ;
      RECT 123.49 212.28 129.98 212.44 ;
      RECT 123.47 215.68 129.98 215.84 ;
      RECT 123.49 219.08 129.98 219.24 ;
      RECT 123.47 222.48 129.98 222.64 ;
      RECT 123.49 225.88 129.98 226.04 ;
      RECT 123.47 229.28 129.98 229.44 ;
      RECT 123.49 232.68 129.98 232.84 ;
      RECT 123.47 236.08 129.98 236.24 ;
      RECT 123.49 239.48 129.98 239.64 ;
      RECT 123.47 242.88 129.98 243.04 ;
      RECT 123.49 246.28 129.98 246.44 ;
      RECT 123.47 249.68 129.98 249.84 ;
      RECT 123.49 253.08 129.98 253.24 ;
      RECT 123.47 256.48 129.98 256.64 ;
      RECT 123.49 259.88 129.98 260.04 ;
      RECT 123.47 263.28 129.98 263.44 ;
      RECT 123.49 266.68 129.98 266.84 ;
      RECT 123.47 270.08 129.98 270.24 ;
      RECT 123.49 273.48 129.98 273.64 ;
      RECT 123.47 276.88 129.98 277.04 ;
      RECT 123.49 280.28 129.98 280.44 ;
      RECT 123.47 283.68 129.98 283.84 ;
      RECT 123.49 287.08 129.98 287.24 ;
      RECT 123.47 290.48 129.98 290.64 ;
      RECT 123.49 293.88 129.98 294.04 ;
      RECT 123.47 297.28 129.98 297.44 ;
      RECT 123.49 300.68 129.98 300.84 ;
      RECT 123.47 304.08 129.98 304.24 ;
      RECT 123.49 307.48 129.98 307.64 ;
      RECT 123.47 310.88 129.98 311.04 ;
      RECT 123.49 314.28 129.98 314.44 ;
      RECT 123.47 317.68 129.98 317.84 ;
      RECT 123.49 321.08 129.98 321.24 ;
      RECT 123.47 324.48 129.98 324.64 ;
      RECT 123.49 327.88 129.98 328.04 ;
      RECT 123.47 331.28 129.98 331.44 ;
      RECT 123.49 334.68 129.98 334.84 ;
      RECT 123.47 338.08 129.98 338.24 ;
      RECT 123.49 341.48 129.98 341.64 ;
      RECT 123.47 344.88 129.98 345.04 ;
      RECT 123.49 348.28 129.98 348.44 ;
      RECT 123.47 351.68 129.98 351.84 ;
      RECT 123.49 355.08 129.98 355.24 ;
      RECT 123.47 358.48 129.98 358.64 ;
      RECT 123.49 361.88 129.98 362.04 ;
      RECT 123.47 365.28 129.98 365.44 ;
      RECT 123.49 368.68 129.98 368.84 ;
      RECT 123.47 372.08 129.98 372.24 ;
      RECT 123.49 375.48 129.98 375.64 ;
      RECT 123.47 378.88 129.98 379.04 ;
      RECT 123.49 382.28 129.98 382.44 ;
      RECT 123.47 385.68 129.98 385.84 ;
      RECT 123.49 389.08 129.98 389.24 ;
      RECT 123.47 392.48 129.98 392.64 ;
      RECT 123.49 395.88 129.98 396.04 ;
      RECT 123.47 399.28 129.98 399.44 ;
      RECT 123.49 402.68 129.98 402.84 ;
      RECT 123.47 406.08 129.98 406.24 ;
      RECT 123.49 409.48 129.98 409.64 ;
      RECT 123.47 412.88 129.98 413.04 ;
      RECT 123.49 416.28 129.98 416.44 ;
      RECT 123.47 419.68 129.98 419.84 ;
      RECT 123.49 423.08 129.98 423.24 ;
      RECT 123.47 426.48 129.98 426.64 ;
      RECT 123.49 429.88 129.98 430.04 ;
      RECT 123.47 433.28 129.98 433.44 ;
      RECT 123.49 436.68 129.98 436.84 ;
      RECT 123.47 440.08 129.98 440.24 ;
      RECT 123.49 443.48 129.98 443.64 ;
      RECT 123.47 446.88 129.98 447.04 ;
      RECT 123.49 450.28 129.98 450.44 ;
      RECT 123.47 453.68 129.98 453.84 ;
      RECT 123.49 457.08 129.98 457.24 ;
      RECT 123.47 460.48 129.98 460.64 ;
      RECT 123.49 463.88 129.98 464.04 ;
      RECT 123.47 467.28 129.98 467.44 ;
      RECT 123.49 470.68 129.98 470.84 ;
      RECT 123.47 474.08 129.98 474.24 ;
      RECT 123.49 477.48 129.98 477.64 ;
      RECT 123.47 480.88 129.98 481.04 ;
      RECT 123.49 484.28 129.98 484.44 ;
      RECT 123.47 487.68 129.98 487.84 ;
      RECT 123.49 491.08 129.98 491.24 ;
      RECT 123.47 494.48 129.98 494.64 ;
      RECT 123.49 497.88 129.98 498.04 ;
      RECT 123.47 501.28 129.98 501.44 ;
      RECT 127.98 505.48 129.95 505.8 ;
      RECT 129.53 12.63 129.69 17.44 ;
      RECT 129.53 17.6 129.69 20.88 ;
      RECT 129.53 32.85 129.69 36.97 ;
      RECT 129.53 40.73 129.69 41.55 ;
      RECT 129.53 60.41 129.69 64 ;
      RECT 127.88 70.38 129.36 70.6 ;
      RECT 127.88 71.92 129.36 72.14 ;
      RECT 127.88 73.78 129.36 74 ;
      RECT 127.88 75.32 129.36 75.54 ;
      RECT 127.88 77.18 129.36 77.4 ;
      RECT 127.88 78.72 129.36 78.94 ;
      RECT 127.88 80.58 129.36 80.8 ;
      RECT 127.88 82.12 129.36 82.34 ;
      RECT 127.88 83.98 129.36 84.2 ;
      RECT 127.88 85.52 129.36 85.74 ;
      RECT 127.88 87.38 129.36 87.6 ;
      RECT 127.88 88.92 129.36 89.14 ;
      RECT 127.88 90.78 129.36 91 ;
      RECT 127.88 92.32 129.36 92.54 ;
      RECT 127.88 94.18 129.36 94.4 ;
      RECT 127.88 95.72 129.36 95.94 ;
      RECT 127.88 97.58 129.36 97.8 ;
      RECT 127.88 99.12 129.36 99.34 ;
      RECT 127.88 100.98 129.36 101.2 ;
      RECT 127.88 102.52 129.36 102.74 ;
      RECT 127.88 104.38 129.36 104.6 ;
      RECT 127.88 105.92 129.36 106.14 ;
      RECT 127.88 107.78 129.36 108 ;
      RECT 127.88 109.32 129.36 109.54 ;
      RECT 127.88 111.18 129.36 111.4 ;
      RECT 127.88 112.72 129.36 112.94 ;
      RECT 127.88 114.58 129.36 114.8 ;
      RECT 127.88 116.12 129.36 116.34 ;
      RECT 127.88 117.98 129.36 118.2 ;
      RECT 127.88 119.52 129.36 119.74 ;
      RECT 127.88 121.38 129.36 121.6 ;
      RECT 127.88 122.92 129.36 123.14 ;
      RECT 127.88 124.78 129.36 125 ;
      RECT 127.88 126.32 129.36 126.54 ;
      RECT 127.88 128.18 129.36 128.4 ;
      RECT 127.88 129.72 129.36 129.94 ;
      RECT 127.88 131.58 129.36 131.8 ;
      RECT 127.88 133.12 129.36 133.34 ;
      RECT 127.88 134.98 129.36 135.2 ;
      RECT 127.88 136.52 129.36 136.74 ;
      RECT 127.88 138.38 129.36 138.6 ;
      RECT 127.88 139.92 129.36 140.14 ;
      RECT 127.88 141.78 129.36 142 ;
      RECT 127.88 143.32 129.36 143.54 ;
      RECT 127.88 145.18 129.36 145.4 ;
      RECT 127.88 146.72 129.36 146.94 ;
      RECT 127.88 148.58 129.36 148.8 ;
      RECT 127.88 150.12 129.36 150.34 ;
      RECT 127.88 151.98 129.36 152.2 ;
      RECT 127.88 153.52 129.36 153.74 ;
      RECT 127.88 155.38 129.36 155.6 ;
      RECT 127.88 156.92 129.36 157.14 ;
      RECT 127.88 158.78 129.36 159 ;
      RECT 127.88 160.32 129.36 160.54 ;
      RECT 127.88 162.18 129.36 162.4 ;
      RECT 127.88 163.72 129.36 163.94 ;
      RECT 127.88 165.58 129.36 165.8 ;
      RECT 127.88 167.12 129.36 167.34 ;
      RECT 127.88 168.98 129.36 169.2 ;
      RECT 127.88 170.52 129.36 170.74 ;
      RECT 127.88 172.38 129.36 172.6 ;
      RECT 127.88 173.92 129.36 174.14 ;
      RECT 127.88 175.78 129.36 176 ;
      RECT 127.88 177.32 129.36 177.54 ;
      RECT 127.88 179.18 129.36 179.4 ;
      RECT 127.88 180.72 129.36 180.94 ;
      RECT 127.88 182.58 129.36 182.8 ;
      RECT 127.88 184.12 129.36 184.34 ;
      RECT 127.88 185.98 129.36 186.2 ;
      RECT 127.88 187.52 129.36 187.74 ;
      RECT 127.88 189.38 129.36 189.6 ;
      RECT 127.88 190.92 129.36 191.14 ;
      RECT 127.88 192.78 129.36 193 ;
      RECT 127.88 194.32 129.36 194.54 ;
      RECT 127.88 196.18 129.36 196.4 ;
      RECT 127.88 197.72 129.36 197.94 ;
      RECT 127.88 199.58 129.36 199.8 ;
      RECT 127.88 201.12 129.36 201.34 ;
      RECT 127.88 202.98 129.36 203.2 ;
      RECT 127.88 204.52 129.36 204.74 ;
      RECT 127.88 206.38 129.36 206.6 ;
      RECT 127.88 207.92 129.36 208.14 ;
      RECT 127.88 209.78 129.36 210 ;
      RECT 127.88 211.32 129.36 211.54 ;
      RECT 127.88 213.18 129.36 213.4 ;
      RECT 127.88 214.72 129.36 214.94 ;
      RECT 127.88 216.58 129.36 216.8 ;
      RECT 127.88 218.12 129.36 218.34 ;
      RECT 127.88 219.98 129.36 220.2 ;
      RECT 127.88 221.52 129.36 221.74 ;
      RECT 127.88 223.38 129.36 223.6 ;
      RECT 127.88 224.92 129.36 225.14 ;
      RECT 127.88 226.78 129.36 227 ;
      RECT 127.88 228.32 129.36 228.54 ;
      RECT 127.88 230.18 129.36 230.4 ;
      RECT 127.88 231.72 129.36 231.94 ;
      RECT 127.88 233.58 129.36 233.8 ;
      RECT 127.88 235.12 129.36 235.34 ;
      RECT 127.88 236.98 129.36 237.2 ;
      RECT 127.88 238.52 129.36 238.74 ;
      RECT 127.88 240.38 129.36 240.6 ;
      RECT 127.88 241.92 129.36 242.14 ;
      RECT 127.88 243.78 129.36 244 ;
      RECT 127.88 245.32 129.36 245.54 ;
      RECT 127.88 247.18 129.36 247.4 ;
      RECT 127.88 248.72 129.36 248.94 ;
      RECT 127.88 250.58 129.36 250.8 ;
      RECT 127.88 252.12 129.36 252.34 ;
      RECT 127.88 253.98 129.36 254.2 ;
      RECT 127.88 255.52 129.36 255.74 ;
      RECT 127.88 257.38 129.36 257.6 ;
      RECT 127.88 258.92 129.36 259.14 ;
      RECT 127.88 260.78 129.36 261 ;
      RECT 127.88 262.32 129.36 262.54 ;
      RECT 127.88 264.18 129.36 264.4 ;
      RECT 127.88 265.72 129.36 265.94 ;
      RECT 127.88 267.58 129.36 267.8 ;
      RECT 127.88 269.12 129.36 269.34 ;
      RECT 127.88 270.98 129.36 271.2 ;
      RECT 127.88 272.52 129.36 272.74 ;
      RECT 127.88 274.38 129.36 274.6 ;
      RECT 127.88 275.92 129.36 276.14 ;
      RECT 127.88 277.78 129.36 278 ;
      RECT 127.88 279.32 129.36 279.54 ;
      RECT 127.88 281.18 129.36 281.4 ;
      RECT 127.88 282.72 129.36 282.94 ;
      RECT 127.88 284.58 129.36 284.8 ;
      RECT 127.88 286.12 129.36 286.34 ;
      RECT 127.88 287.98 129.36 288.2 ;
      RECT 127.88 289.52 129.36 289.74 ;
      RECT 127.88 291.38 129.36 291.6 ;
      RECT 127.88 292.92 129.36 293.14 ;
      RECT 127.88 294.78 129.36 295 ;
      RECT 127.88 296.32 129.36 296.54 ;
      RECT 127.88 298.18 129.36 298.4 ;
      RECT 127.88 299.72 129.36 299.94 ;
      RECT 127.88 301.58 129.36 301.8 ;
      RECT 127.88 303.12 129.36 303.34 ;
      RECT 127.88 304.98 129.36 305.2 ;
      RECT 127.88 306.52 129.36 306.74 ;
      RECT 127.88 308.38 129.36 308.6 ;
      RECT 127.88 309.92 129.36 310.14 ;
      RECT 127.88 311.78 129.36 312 ;
      RECT 127.88 313.32 129.36 313.54 ;
      RECT 127.88 315.18 129.36 315.4 ;
      RECT 127.88 316.72 129.36 316.94 ;
      RECT 127.88 318.58 129.36 318.8 ;
      RECT 127.88 320.12 129.36 320.34 ;
      RECT 127.88 321.98 129.36 322.2 ;
      RECT 127.88 323.52 129.36 323.74 ;
      RECT 127.88 325.38 129.36 325.6 ;
      RECT 127.88 326.92 129.36 327.14 ;
      RECT 127.88 328.78 129.36 329 ;
      RECT 127.88 330.32 129.36 330.54 ;
      RECT 127.88 332.18 129.36 332.4 ;
      RECT 127.88 333.72 129.36 333.94 ;
      RECT 127.88 335.58 129.36 335.8 ;
      RECT 127.88 337.12 129.36 337.34 ;
      RECT 127.88 338.98 129.36 339.2 ;
      RECT 127.88 340.52 129.36 340.74 ;
      RECT 127.88 342.38 129.36 342.6 ;
      RECT 127.88 343.92 129.36 344.14 ;
      RECT 127.88 345.78 129.36 346 ;
      RECT 127.88 347.32 129.36 347.54 ;
      RECT 127.88 349.18 129.36 349.4 ;
      RECT 127.88 350.72 129.36 350.94 ;
      RECT 127.88 352.58 129.36 352.8 ;
      RECT 127.88 354.12 129.36 354.34 ;
      RECT 127.88 355.98 129.36 356.2 ;
      RECT 127.88 357.52 129.36 357.74 ;
      RECT 127.88 359.38 129.36 359.6 ;
      RECT 127.88 360.92 129.36 361.14 ;
      RECT 127.88 362.78 129.36 363 ;
      RECT 127.88 364.32 129.36 364.54 ;
      RECT 127.88 366.18 129.36 366.4 ;
      RECT 127.88 367.72 129.36 367.94 ;
      RECT 127.88 369.58 129.36 369.8 ;
      RECT 127.88 371.12 129.36 371.34 ;
      RECT 127.88 372.98 129.36 373.2 ;
      RECT 127.88 374.52 129.36 374.74 ;
      RECT 127.88 376.38 129.36 376.6 ;
      RECT 127.88 377.92 129.36 378.14 ;
      RECT 127.88 379.78 129.36 380 ;
      RECT 127.88 381.32 129.36 381.54 ;
      RECT 127.88 383.18 129.36 383.4 ;
      RECT 127.88 384.72 129.36 384.94 ;
      RECT 127.88 386.58 129.36 386.8 ;
      RECT 127.88 388.12 129.36 388.34 ;
      RECT 127.88 389.98 129.36 390.2 ;
      RECT 127.88 391.52 129.36 391.74 ;
      RECT 127.88 393.38 129.36 393.6 ;
      RECT 127.88 394.92 129.36 395.14 ;
      RECT 127.88 396.78 129.36 397 ;
      RECT 127.88 398.32 129.36 398.54 ;
      RECT 127.88 400.18 129.36 400.4 ;
      RECT 127.88 401.72 129.36 401.94 ;
      RECT 127.88 403.58 129.36 403.8 ;
      RECT 127.88 405.12 129.36 405.34 ;
      RECT 127.88 406.98 129.36 407.2 ;
      RECT 127.88 408.52 129.36 408.74 ;
      RECT 127.88 410.38 129.36 410.6 ;
      RECT 127.88 411.92 129.36 412.14 ;
      RECT 127.88 413.78 129.36 414 ;
      RECT 127.88 415.32 129.36 415.54 ;
      RECT 127.88 417.18 129.36 417.4 ;
      RECT 127.88 418.72 129.36 418.94 ;
      RECT 127.88 420.58 129.36 420.8 ;
      RECT 127.88 422.12 129.36 422.34 ;
      RECT 127.88 423.98 129.36 424.2 ;
      RECT 127.88 425.52 129.36 425.74 ;
      RECT 127.88 427.38 129.36 427.6 ;
      RECT 127.88 428.92 129.36 429.14 ;
      RECT 127.88 430.78 129.36 431 ;
      RECT 127.88 432.32 129.36 432.54 ;
      RECT 127.88 434.18 129.36 434.4 ;
      RECT 127.88 435.72 129.36 435.94 ;
      RECT 127.88 437.58 129.36 437.8 ;
      RECT 127.88 439.12 129.36 439.34 ;
      RECT 127.88 440.98 129.36 441.2 ;
      RECT 127.88 442.52 129.36 442.74 ;
      RECT 127.88 444.38 129.36 444.6 ;
      RECT 127.88 445.92 129.36 446.14 ;
      RECT 127.88 447.78 129.36 448 ;
      RECT 127.88 449.32 129.36 449.54 ;
      RECT 127.88 451.18 129.36 451.4 ;
      RECT 127.88 452.72 129.36 452.94 ;
      RECT 127.88 454.58 129.36 454.8 ;
      RECT 127.88 456.12 129.36 456.34 ;
      RECT 127.88 457.98 129.36 458.2 ;
      RECT 127.88 459.52 129.36 459.74 ;
      RECT 127.88 461.38 129.36 461.6 ;
      RECT 127.88 462.92 129.36 463.14 ;
      RECT 127.88 464.78 129.36 465 ;
      RECT 127.88 466.32 129.36 466.54 ;
      RECT 127.88 468.18 129.36 468.4 ;
      RECT 127.88 469.72 129.36 469.94 ;
      RECT 127.88 471.58 129.36 471.8 ;
      RECT 127.88 473.12 129.36 473.34 ;
      RECT 127.88 474.98 129.36 475.2 ;
      RECT 127.88 476.52 129.36 476.74 ;
      RECT 127.88 478.38 129.36 478.6 ;
      RECT 127.88 479.92 129.36 480.14 ;
      RECT 127.88 481.78 129.36 482 ;
      RECT 127.88 483.32 129.36 483.54 ;
      RECT 127.88 485.18 129.36 485.4 ;
      RECT 127.88 486.72 129.36 486.94 ;
      RECT 127.88 488.58 129.36 488.8 ;
      RECT 127.88 490.12 129.36 490.34 ;
      RECT 127.88 491.98 129.36 492.2 ;
      RECT 127.88 493.52 129.36 493.74 ;
      RECT 127.88 495.38 129.36 495.6 ;
      RECT 127.88 496.92 129.36 497.14 ;
      RECT 127.88 498.78 129.36 499 ;
      RECT 127.88 500.32 129.36 500.54 ;
      RECT 127.88 502.18 129.36 502.4 ;
      RECT 127.88 503.72 129.36 503.94 ;
      RECT 129.05 9.61 129.21 14.44 ;
      RECT 128.84 37.58 129.03 38.41 ;
      RECT 128.71 38.57 128.87 40.5 ;
      RECT 128.42 37.58 128.59 38.41 ;
      RECT 128.31 17.46 128.47 20.88 ;
      RECT 128.31 61.17 128.47 64.59 ;
      RECT 127.57 23.99 128.25 24.21 ;
      RECT 127.57 57.84 128.25 58.06 ;
      RECT 127.74 7.04 128.06 7.36 ;
      RECT 124.81 510.54 127.61 510.94 ;
      RECT 127.24 37.58 127.52 38.41 ;
      RECT 127.35 17.46 127.51 20.88 ;
      RECT 127.35 61.17 127.51 64.59 ;
      RECT 125.21 6.24 127.19 6.84 ;
      RECT 126.95 38.57 127.11 40.5 ;
      RECT 126.79 37.58 127.08 38.41 ;
      RECT 126.87 30.54 127.03 32.2 ;
      RECT 126.87 50.09 127.03 51.7 ;
      RECT 126.61 9.61 126.77 14.44 ;
      RECT 126.1 23.97 126.32 24.48 ;
      RECT 126.1 57.58 126.32 58.08 ;
      RECT 126.13 12.63 126.29 17.44 ;
      RECT 126.13 31.09 126.29 36.97 ;
      RECT 126.13 40.73 126.29 41.55 ;
      RECT 126.13 45.65 126.29 51.3 ;
      RECT 125.34 37.58 125.63 38.41 ;
      RECT 125.39 30.54 125.55 32.2 ;
      RECT 125.39 50.09 125.55 51.7 ;
      RECT 125.31 38.57 125.47 40.5 ;
      RECT 124.9 37.58 125.18 38.41 ;
      RECT 124.91 14.52 125.07 16.86 ;
      RECT 124.91 17.46 125.07 20.88 ;
      RECT 124.91 61.17 125.07 64.59 ;
      RECT 124.17 23.99 124.85 24.21 ;
      RECT 124.17 57.84 124.85 58.06 ;
      RECT 121.24 71.18 124.14 71.34 ;
      RECT 121.24 74.58 124.14 74.74 ;
      RECT 121.24 77.98 124.14 78.14 ;
      RECT 121.24 81.38 124.14 81.54 ;
      RECT 121.24 84.78 124.14 84.94 ;
      RECT 121.24 88.18 124.14 88.34 ;
      RECT 121.24 91.58 124.14 91.74 ;
      RECT 121.24 94.98 124.14 95.14 ;
      RECT 121.24 98.38 124.14 98.54 ;
      RECT 121.24 101.78 124.14 101.94 ;
      RECT 121.24 105.18 124.14 105.34 ;
      RECT 121.24 108.58 124.14 108.74 ;
      RECT 121.24 111.98 124.14 112.14 ;
      RECT 121.24 115.38 124.14 115.54 ;
      RECT 121.24 118.78 124.14 118.94 ;
      RECT 121.24 122.18 124.14 122.34 ;
      RECT 121.24 125.58 124.14 125.74 ;
      RECT 121.24 128.98 124.14 129.14 ;
      RECT 121.24 132.38 124.14 132.54 ;
      RECT 121.24 135.78 124.14 135.94 ;
      RECT 121.24 139.18 124.14 139.34 ;
      RECT 121.24 142.58 124.14 142.74 ;
      RECT 121.24 145.98 124.14 146.14 ;
      RECT 121.24 149.38 124.14 149.54 ;
      RECT 121.24 152.78 124.14 152.94 ;
      RECT 121.24 156.18 124.14 156.34 ;
      RECT 121.24 159.58 124.14 159.74 ;
      RECT 121.24 162.98 124.14 163.14 ;
      RECT 121.24 166.38 124.14 166.54 ;
      RECT 121.24 169.78 124.14 169.94 ;
      RECT 121.24 173.18 124.14 173.34 ;
      RECT 121.24 176.58 124.14 176.74 ;
      RECT 121.24 179.98 124.14 180.14 ;
      RECT 121.24 183.38 124.14 183.54 ;
      RECT 121.24 186.78 124.14 186.94 ;
      RECT 121.24 190.18 124.14 190.34 ;
      RECT 121.24 193.58 124.14 193.74 ;
      RECT 121.24 196.98 124.14 197.14 ;
      RECT 121.24 200.38 124.14 200.54 ;
      RECT 121.24 203.78 124.14 203.94 ;
      RECT 121.24 207.18 124.14 207.34 ;
      RECT 121.24 210.58 124.14 210.74 ;
      RECT 121.24 213.98 124.14 214.14 ;
      RECT 121.24 217.38 124.14 217.54 ;
      RECT 121.24 220.78 124.14 220.94 ;
      RECT 121.24 224.18 124.14 224.34 ;
      RECT 121.24 227.58 124.14 227.74 ;
      RECT 121.24 230.98 124.14 231.14 ;
      RECT 121.24 234.38 124.14 234.54 ;
      RECT 121.24 237.78 124.14 237.94 ;
      RECT 121.24 241.18 124.14 241.34 ;
      RECT 121.24 244.58 124.14 244.74 ;
      RECT 121.24 247.98 124.14 248.14 ;
      RECT 121.24 251.38 124.14 251.54 ;
      RECT 121.24 254.78 124.14 254.94 ;
      RECT 121.24 258.18 124.14 258.34 ;
      RECT 121.24 261.58 124.14 261.74 ;
      RECT 121.24 264.98 124.14 265.14 ;
      RECT 121.24 268.38 124.14 268.54 ;
      RECT 121.24 271.78 124.14 271.94 ;
      RECT 121.24 275.18 124.14 275.34 ;
      RECT 121.24 278.58 124.14 278.74 ;
      RECT 121.24 281.98 124.14 282.14 ;
      RECT 121.24 285.38 124.14 285.54 ;
      RECT 121.24 288.78 124.14 288.94 ;
      RECT 121.24 292.18 124.14 292.34 ;
      RECT 121.24 295.58 124.14 295.74 ;
      RECT 121.24 298.98 124.14 299.14 ;
      RECT 121.24 302.38 124.14 302.54 ;
      RECT 121.24 305.78 124.14 305.94 ;
      RECT 121.24 309.18 124.14 309.34 ;
      RECT 121.24 312.58 124.14 312.74 ;
      RECT 121.24 315.98 124.14 316.14 ;
      RECT 121.24 319.38 124.14 319.54 ;
      RECT 121.24 322.78 124.14 322.94 ;
      RECT 121.24 326.18 124.14 326.34 ;
      RECT 121.24 329.58 124.14 329.74 ;
      RECT 121.24 332.98 124.14 333.14 ;
      RECT 121.24 336.38 124.14 336.54 ;
      RECT 121.24 339.78 124.14 339.94 ;
      RECT 121.24 343.18 124.14 343.34 ;
      RECT 121.24 346.58 124.14 346.74 ;
      RECT 121.24 349.98 124.14 350.14 ;
      RECT 121.24 353.38 124.14 353.54 ;
      RECT 121.24 356.78 124.14 356.94 ;
      RECT 121.24 360.18 124.14 360.34 ;
      RECT 121.24 363.58 124.14 363.74 ;
      RECT 121.24 366.98 124.14 367.14 ;
      RECT 121.24 370.38 124.14 370.54 ;
      RECT 121.24 373.78 124.14 373.94 ;
      RECT 121.24 377.18 124.14 377.34 ;
      RECT 121.24 380.58 124.14 380.74 ;
      RECT 121.24 383.98 124.14 384.14 ;
      RECT 121.24 387.38 124.14 387.54 ;
      RECT 121.24 390.78 124.14 390.94 ;
      RECT 121.24 394.18 124.14 394.34 ;
      RECT 121.24 397.58 124.14 397.74 ;
      RECT 121.24 400.98 124.14 401.14 ;
      RECT 121.24 404.38 124.14 404.54 ;
      RECT 121.24 407.78 124.14 407.94 ;
      RECT 121.24 411.18 124.14 411.34 ;
      RECT 121.24 414.58 124.14 414.74 ;
      RECT 121.24 417.98 124.14 418.14 ;
      RECT 121.24 421.38 124.14 421.54 ;
      RECT 121.24 424.78 124.14 424.94 ;
      RECT 121.24 428.18 124.14 428.34 ;
      RECT 121.24 431.58 124.14 431.74 ;
      RECT 121.24 434.98 124.14 435.14 ;
      RECT 121.24 438.38 124.14 438.54 ;
      RECT 121.24 441.78 124.14 441.94 ;
      RECT 121.24 445.18 124.14 445.34 ;
      RECT 121.24 448.58 124.14 448.74 ;
      RECT 121.24 451.98 124.14 452.14 ;
      RECT 121.24 455.38 124.14 455.54 ;
      RECT 121.24 458.78 124.14 458.94 ;
      RECT 121.24 462.18 124.14 462.34 ;
      RECT 121.24 465.58 124.14 465.74 ;
      RECT 121.24 468.98 124.14 469.14 ;
      RECT 121.24 472.38 124.14 472.54 ;
      RECT 121.24 475.78 124.14 475.94 ;
      RECT 121.24 479.18 124.14 479.34 ;
      RECT 121.24 482.58 124.14 482.74 ;
      RECT 121.24 485.98 124.14 486.14 ;
      RECT 121.24 489.38 124.14 489.54 ;
      RECT 121.24 492.78 124.14 492.94 ;
      RECT 121.24 496.18 124.14 496.34 ;
      RECT 121.24 499.58 124.14 499.74 ;
      RECT 121.24 502.98 124.14 503.14 ;
      RECT 123.95 14.52 124.11 16.86 ;
      RECT 123.95 17.46 124.11 20.88 ;
      RECT 123.95 61.17 124.11 64.59 ;
      RECT 123.83 37.58 124 38.41 ;
      RECT 121.83 6.24 123.81 6.84 ;
      RECT 123.55 38.57 123.71 40.5 ;
      RECT 123.39 37.58 123.58 38.41 ;
      RECT 122.73 12.63 122.89 17.44 ;
      RECT 122.73 17.6 122.89 20.88 ;
      RECT 122.73 32.85 122.89 36.97 ;
      RECT 122.73 40.73 122.89 41.55 ;
      RECT 122.73 60.41 122.89 64 ;
      RECT 122.25 9.61 122.41 14.44 ;
      RECT 122.04 37.58 122.23 38.41 ;
      RECT 121.91 38.57 122.07 40.5 ;
      RECT 121.62 37.58 121.79 38.41 ;
      RECT 121.51 17.46 121.67 20.88 ;
      RECT 121.51 61.17 121.67 64.59 ;
      RECT 120.77 23.99 121.45 24.21 ;
      RECT 120.77 57.84 121.45 58.06 ;
      RECT 114.94 506.76 121.44 506.92 ;
      RECT 114.94 507.24 121.44 507.4 ;
      RECT 120.94 7.04 121.26 7.36 ;
      RECT 118.01 510.54 120.81 510.94 ;
      RECT 120.44 37.58 120.72 38.41 ;
      RECT 120.55 17.46 120.71 20.88 ;
      RECT 120.55 61.17 120.71 64.59 ;
      RECT 118.43 6.24 120.39 6.84 ;
      RECT 120.15 38.57 120.31 40.5 ;
      RECT 119.99 37.58 120.28 38.41 ;
      RECT 120.07 30.54 120.23 32.2 ;
      RECT 120.07 50.09 120.23 51.7 ;
      RECT 119.81 9.61 119.97 14.44 ;
      RECT 119.3 23.97 119.52 24.48 ;
      RECT 119.3 57.58 119.52 58.08 ;
      RECT 119.33 12.63 119.49 17.44 ;
      RECT 119.33 31.09 119.49 36.97 ;
      RECT 119.33 40.73 119.49 41.55 ;
      RECT 119.33 45.65 119.49 51.3 ;
      RECT 118.85 9.61 119.01 14.44 ;
      RECT 117.82 71.23 118.92 71.39 ;
      RECT 117.82 74.53 118.92 74.69 ;
      RECT 117.82 78.03 118.92 78.19 ;
      RECT 117.82 81.33 118.92 81.49 ;
      RECT 117.82 84.83 118.92 84.99 ;
      RECT 117.82 88.13 118.92 88.29 ;
      RECT 117.82 91.63 118.92 91.79 ;
      RECT 117.82 94.93 118.92 95.09 ;
      RECT 117.82 98.43 118.92 98.59 ;
      RECT 117.82 101.73 118.92 101.89 ;
      RECT 117.82 105.23 118.92 105.39 ;
      RECT 117.82 108.53 118.92 108.69 ;
      RECT 117.82 112.03 118.92 112.19 ;
      RECT 117.82 115.33 118.92 115.49 ;
      RECT 117.82 118.83 118.92 118.99 ;
      RECT 117.82 122.13 118.92 122.29 ;
      RECT 117.82 125.63 118.92 125.79 ;
      RECT 117.82 128.93 118.92 129.09 ;
      RECT 117.82 132.43 118.92 132.59 ;
      RECT 117.82 135.73 118.92 135.89 ;
      RECT 117.82 139.23 118.92 139.39 ;
      RECT 117.82 142.53 118.92 142.69 ;
      RECT 117.82 146.03 118.92 146.19 ;
      RECT 117.82 149.33 118.92 149.49 ;
      RECT 117.82 152.83 118.92 152.99 ;
      RECT 117.82 156.13 118.92 156.29 ;
      RECT 117.82 159.63 118.92 159.79 ;
      RECT 117.82 162.93 118.92 163.09 ;
      RECT 117.82 166.43 118.92 166.59 ;
      RECT 117.82 169.73 118.92 169.89 ;
      RECT 117.82 173.23 118.92 173.39 ;
      RECT 117.82 176.53 118.92 176.69 ;
      RECT 117.82 180.03 118.92 180.19 ;
      RECT 117.82 183.33 118.92 183.49 ;
      RECT 117.82 186.83 118.92 186.99 ;
      RECT 117.82 190.13 118.92 190.29 ;
      RECT 117.82 193.63 118.92 193.79 ;
      RECT 117.82 196.93 118.92 197.09 ;
      RECT 117.82 200.43 118.92 200.59 ;
      RECT 117.82 203.73 118.92 203.89 ;
      RECT 117.82 207.23 118.92 207.39 ;
      RECT 117.82 210.53 118.92 210.69 ;
      RECT 117.82 214.03 118.92 214.19 ;
      RECT 117.82 217.33 118.92 217.49 ;
      RECT 117.82 220.83 118.92 220.99 ;
      RECT 117.82 224.13 118.92 224.29 ;
      RECT 117.82 227.63 118.92 227.79 ;
      RECT 117.82 230.93 118.92 231.09 ;
      RECT 117.82 234.43 118.92 234.59 ;
      RECT 117.82 237.73 118.92 237.89 ;
      RECT 117.82 241.23 118.92 241.39 ;
      RECT 117.82 244.53 118.92 244.69 ;
      RECT 117.82 248.03 118.92 248.19 ;
      RECT 117.82 251.33 118.92 251.49 ;
      RECT 117.82 254.83 118.92 254.99 ;
      RECT 117.82 258.13 118.92 258.29 ;
      RECT 117.82 261.63 118.92 261.79 ;
      RECT 117.82 264.93 118.92 265.09 ;
      RECT 117.82 268.43 118.92 268.59 ;
      RECT 117.82 271.73 118.92 271.89 ;
      RECT 117.82 275.23 118.92 275.39 ;
      RECT 117.82 278.53 118.92 278.69 ;
      RECT 117.82 282.03 118.92 282.19 ;
      RECT 117.82 285.33 118.92 285.49 ;
      RECT 117.82 288.83 118.92 288.99 ;
      RECT 117.82 292.13 118.92 292.29 ;
      RECT 117.82 295.63 118.92 295.79 ;
      RECT 117.82 298.93 118.92 299.09 ;
      RECT 117.82 302.43 118.92 302.59 ;
      RECT 117.82 305.73 118.92 305.89 ;
      RECT 117.82 309.23 118.92 309.39 ;
      RECT 117.82 312.53 118.92 312.69 ;
      RECT 117.82 316.03 118.92 316.19 ;
      RECT 117.82 319.33 118.92 319.49 ;
      RECT 117.82 322.83 118.92 322.99 ;
      RECT 117.82 326.13 118.92 326.29 ;
      RECT 117.82 329.63 118.92 329.79 ;
      RECT 117.82 332.93 118.92 333.09 ;
      RECT 117.82 336.43 118.92 336.59 ;
      RECT 117.82 339.73 118.92 339.89 ;
      RECT 117.82 343.23 118.92 343.39 ;
      RECT 117.82 346.53 118.92 346.69 ;
      RECT 117.82 350.03 118.92 350.19 ;
      RECT 117.82 353.33 118.92 353.49 ;
      RECT 117.82 356.83 118.92 356.99 ;
      RECT 117.82 360.13 118.92 360.29 ;
      RECT 117.82 363.63 118.92 363.79 ;
      RECT 117.82 366.93 118.92 367.09 ;
      RECT 117.82 370.43 118.92 370.59 ;
      RECT 117.82 373.73 118.92 373.89 ;
      RECT 117.82 377.23 118.92 377.39 ;
      RECT 117.82 380.53 118.92 380.69 ;
      RECT 117.82 384.03 118.92 384.19 ;
      RECT 117.82 387.33 118.92 387.49 ;
      RECT 117.82 390.83 118.92 390.99 ;
      RECT 117.82 394.13 118.92 394.29 ;
      RECT 117.82 397.63 118.92 397.79 ;
      RECT 117.82 400.93 118.92 401.09 ;
      RECT 117.82 404.43 118.92 404.59 ;
      RECT 117.82 407.73 118.92 407.89 ;
      RECT 117.82 411.23 118.92 411.39 ;
      RECT 117.82 414.53 118.92 414.69 ;
      RECT 117.82 418.03 118.92 418.19 ;
      RECT 117.82 421.33 118.92 421.49 ;
      RECT 117.82 424.83 118.92 424.99 ;
      RECT 117.82 428.13 118.92 428.29 ;
      RECT 117.82 431.63 118.92 431.79 ;
      RECT 117.82 434.93 118.92 435.09 ;
      RECT 117.82 438.43 118.92 438.59 ;
      RECT 117.82 441.73 118.92 441.89 ;
      RECT 117.82 445.23 118.92 445.39 ;
      RECT 117.82 448.53 118.92 448.69 ;
      RECT 117.82 452.03 118.92 452.19 ;
      RECT 117.82 455.33 118.92 455.49 ;
      RECT 117.82 458.83 118.92 458.99 ;
      RECT 117.82 462.13 118.92 462.29 ;
      RECT 117.82 465.63 118.92 465.79 ;
      RECT 117.82 468.93 118.92 469.09 ;
      RECT 117.82 472.43 118.92 472.59 ;
      RECT 117.82 475.73 118.92 475.89 ;
      RECT 117.82 479.23 118.92 479.39 ;
      RECT 117.82 482.53 118.92 482.69 ;
      RECT 117.82 486.03 118.92 486.19 ;
      RECT 117.82 489.33 118.92 489.49 ;
      RECT 117.82 492.83 118.92 492.99 ;
      RECT 117.82 496.13 118.92 496.29 ;
      RECT 117.82 499.63 118.92 499.79 ;
      RECT 117.82 502.93 118.92 503.09 ;
      RECT 118.54 37.58 118.83 38.41 ;
      RECT 118.59 30.54 118.75 32.2 ;
      RECT 118.59 50.09 118.75 51.7 ;
      RECT 118.51 38.57 118.67 40.5 ;
      RECT 118.1 37.58 118.38 38.41 ;
      RECT 118.11 17.46 118.27 20.88 ;
      RECT 118.11 61.17 118.27 64.59 ;
      RECT 117.37 23.99 118.05 24.21 ;
      RECT 117.37 57.84 118.05 58.06 ;
      RECT 117.56 7.04 117.88 7.36 ;
      RECT 116.41 71.23 117.66 71.39 ;
      RECT 116.41 74.53 117.66 74.69 ;
      RECT 116.41 78.03 117.66 78.19 ;
      RECT 116.41 81.33 117.66 81.49 ;
      RECT 116.41 84.83 117.66 84.99 ;
      RECT 116.41 88.13 117.66 88.29 ;
      RECT 116.41 91.63 117.66 91.79 ;
      RECT 116.41 94.93 117.66 95.09 ;
      RECT 116.41 98.43 117.66 98.59 ;
      RECT 116.41 101.73 117.66 101.89 ;
      RECT 116.41 105.23 117.66 105.39 ;
      RECT 116.41 108.53 117.66 108.69 ;
      RECT 116.41 112.03 117.66 112.19 ;
      RECT 116.41 115.33 117.66 115.49 ;
      RECT 116.41 118.83 117.66 118.99 ;
      RECT 116.41 122.13 117.66 122.29 ;
      RECT 116.41 125.63 117.66 125.79 ;
      RECT 116.41 128.93 117.66 129.09 ;
      RECT 116.41 132.43 117.66 132.59 ;
      RECT 116.41 135.73 117.66 135.89 ;
      RECT 116.41 139.23 117.66 139.39 ;
      RECT 116.41 142.53 117.66 142.69 ;
      RECT 116.41 146.03 117.66 146.19 ;
      RECT 116.41 149.33 117.66 149.49 ;
      RECT 116.41 152.83 117.66 152.99 ;
      RECT 116.41 156.13 117.66 156.29 ;
      RECT 116.41 159.63 117.66 159.79 ;
      RECT 116.41 162.93 117.66 163.09 ;
      RECT 116.41 166.43 117.66 166.59 ;
      RECT 116.41 169.73 117.66 169.89 ;
      RECT 116.41 173.23 117.66 173.39 ;
      RECT 116.41 176.53 117.66 176.69 ;
      RECT 116.41 180.03 117.66 180.19 ;
      RECT 116.41 183.33 117.66 183.49 ;
      RECT 116.41 186.83 117.66 186.99 ;
      RECT 116.41 190.13 117.66 190.29 ;
      RECT 116.41 193.63 117.66 193.79 ;
      RECT 116.41 196.93 117.66 197.09 ;
      RECT 116.41 200.43 117.66 200.59 ;
      RECT 116.41 203.73 117.66 203.89 ;
      RECT 116.41 207.23 117.66 207.39 ;
      RECT 116.41 210.53 117.66 210.69 ;
      RECT 116.41 214.03 117.66 214.19 ;
      RECT 116.41 217.33 117.66 217.49 ;
      RECT 116.41 220.83 117.66 220.99 ;
      RECT 116.41 224.13 117.66 224.29 ;
      RECT 116.41 227.63 117.66 227.79 ;
      RECT 116.41 230.93 117.66 231.09 ;
      RECT 116.41 234.43 117.66 234.59 ;
      RECT 116.41 237.73 117.66 237.89 ;
      RECT 116.41 241.23 117.66 241.39 ;
      RECT 116.41 244.53 117.66 244.69 ;
      RECT 116.41 248.03 117.66 248.19 ;
      RECT 116.41 251.33 117.66 251.49 ;
      RECT 116.41 254.83 117.66 254.99 ;
      RECT 116.41 258.13 117.66 258.29 ;
      RECT 116.41 261.63 117.66 261.79 ;
      RECT 116.41 264.93 117.66 265.09 ;
      RECT 116.41 268.43 117.66 268.59 ;
      RECT 116.41 271.73 117.66 271.89 ;
      RECT 116.41 275.23 117.66 275.39 ;
      RECT 116.41 278.53 117.66 278.69 ;
      RECT 116.41 282.03 117.66 282.19 ;
      RECT 116.41 285.33 117.66 285.49 ;
      RECT 116.41 288.83 117.66 288.99 ;
      RECT 116.41 292.13 117.66 292.29 ;
      RECT 116.41 295.63 117.66 295.79 ;
      RECT 116.41 298.93 117.66 299.09 ;
      RECT 116.41 302.43 117.66 302.59 ;
      RECT 116.41 305.73 117.66 305.89 ;
      RECT 116.41 309.23 117.66 309.39 ;
      RECT 116.41 312.53 117.66 312.69 ;
      RECT 116.41 316.03 117.66 316.19 ;
      RECT 116.41 319.33 117.66 319.49 ;
      RECT 116.41 322.83 117.66 322.99 ;
      RECT 116.41 326.13 117.66 326.29 ;
      RECT 116.41 329.63 117.66 329.79 ;
      RECT 116.41 332.93 117.66 333.09 ;
      RECT 116.41 336.43 117.66 336.59 ;
      RECT 116.41 339.73 117.66 339.89 ;
      RECT 116.41 343.23 117.66 343.39 ;
      RECT 116.41 346.53 117.66 346.69 ;
      RECT 116.41 350.03 117.66 350.19 ;
      RECT 116.41 353.33 117.66 353.49 ;
      RECT 116.41 356.83 117.66 356.99 ;
      RECT 116.41 360.13 117.66 360.29 ;
      RECT 116.41 363.63 117.66 363.79 ;
      RECT 116.41 366.93 117.66 367.09 ;
      RECT 116.41 370.43 117.66 370.59 ;
      RECT 116.41 373.73 117.66 373.89 ;
      RECT 116.41 377.23 117.66 377.39 ;
      RECT 116.41 380.53 117.66 380.69 ;
      RECT 116.41 384.03 117.66 384.19 ;
      RECT 116.41 387.33 117.66 387.49 ;
      RECT 116.41 390.83 117.66 390.99 ;
      RECT 116.41 394.13 117.66 394.29 ;
      RECT 116.41 397.63 117.66 397.79 ;
      RECT 116.41 400.93 117.66 401.09 ;
      RECT 116.41 404.43 117.66 404.59 ;
      RECT 116.41 407.73 117.66 407.89 ;
      RECT 116.41 411.23 117.66 411.39 ;
      RECT 116.41 414.53 117.66 414.69 ;
      RECT 116.41 418.03 117.66 418.19 ;
      RECT 116.41 421.33 117.66 421.49 ;
      RECT 116.41 424.83 117.66 424.99 ;
      RECT 116.41 428.13 117.66 428.29 ;
      RECT 116.41 431.63 117.66 431.79 ;
      RECT 116.41 434.93 117.66 435.09 ;
      RECT 116.41 438.43 117.66 438.59 ;
      RECT 116.41 441.73 117.66 441.89 ;
      RECT 116.41 445.23 117.66 445.39 ;
      RECT 116.41 448.53 117.66 448.69 ;
      RECT 116.41 452.03 117.66 452.19 ;
      RECT 116.41 455.33 117.66 455.49 ;
      RECT 116.41 458.83 117.66 458.99 ;
      RECT 116.41 462.13 117.66 462.29 ;
      RECT 116.41 465.63 117.66 465.79 ;
      RECT 116.41 468.93 117.66 469.09 ;
      RECT 116.41 472.43 117.66 472.59 ;
      RECT 116.41 475.73 117.66 475.89 ;
      RECT 116.41 479.23 117.66 479.39 ;
      RECT 116.41 482.53 117.66 482.69 ;
      RECT 116.41 486.03 117.66 486.19 ;
      RECT 116.41 489.33 117.66 489.49 ;
      RECT 116.41 492.83 117.66 492.99 ;
      RECT 116.41 496.13 117.66 496.29 ;
      RECT 116.41 499.63 117.66 499.79 ;
      RECT 116.76 502.93 117.66 503.09 ;
      RECT 117.15 17.46 117.31 20.88 ;
      RECT 117.15 61.17 117.31 64.59 ;
      RECT 117.03 37.58 117.2 38.41 ;
      RECT 115.03 6.24 116.99 6.84 ;
      RECT 116.75 38.57 116.91 40.5 ;
      RECT 116.59 37.58 116.78 38.41 ;
      RECT 116.41 69.48 116.76 69.64 ;
      RECT 116.41 72.88 116.76 73.04 ;
      RECT 116.41 76.28 116.76 76.44 ;
      RECT 116.41 79.68 116.76 79.84 ;
      RECT 116.41 83.08 116.76 83.24 ;
      RECT 116.41 86.48 116.76 86.64 ;
      RECT 116.41 89.88 116.76 90.04 ;
      RECT 116.41 93.28 116.76 93.44 ;
      RECT 116.41 96.68 116.76 96.84 ;
      RECT 116.41 100.08 116.76 100.24 ;
      RECT 116.41 103.48 116.76 103.64 ;
      RECT 116.41 106.88 116.76 107.04 ;
      RECT 116.41 110.28 116.76 110.44 ;
      RECT 116.41 113.68 116.76 113.84 ;
      RECT 116.41 117.08 116.76 117.24 ;
      RECT 116.41 120.48 116.76 120.64 ;
      RECT 116.41 123.88 116.76 124.04 ;
      RECT 116.41 127.28 116.76 127.44 ;
      RECT 116.41 130.68 116.76 130.84 ;
      RECT 116.41 134.08 116.76 134.24 ;
      RECT 116.41 137.48 116.76 137.64 ;
      RECT 116.41 140.88 116.76 141.04 ;
      RECT 116.41 144.28 116.76 144.44 ;
      RECT 116.41 147.68 116.76 147.84 ;
      RECT 116.41 151.08 116.76 151.24 ;
      RECT 116.41 154.48 116.76 154.64 ;
      RECT 116.41 157.88 116.76 158.04 ;
      RECT 116.41 161.28 116.76 161.44 ;
      RECT 116.41 164.68 116.76 164.84 ;
      RECT 116.41 168.08 116.76 168.24 ;
      RECT 116.41 171.48 116.76 171.64 ;
      RECT 116.41 174.88 116.76 175.04 ;
      RECT 116.41 178.28 116.76 178.44 ;
      RECT 116.41 181.68 116.76 181.84 ;
      RECT 116.41 185.08 116.76 185.24 ;
      RECT 116.41 188.48 116.76 188.64 ;
      RECT 116.41 191.88 116.76 192.04 ;
      RECT 116.41 195.28 116.76 195.44 ;
      RECT 116.41 198.68 116.76 198.84 ;
      RECT 116.41 202.08 116.76 202.24 ;
      RECT 116.41 205.48 116.76 205.64 ;
      RECT 116.41 208.88 116.76 209.04 ;
      RECT 116.41 212.28 116.76 212.44 ;
      RECT 116.41 215.68 116.76 215.84 ;
      RECT 116.41 219.08 116.76 219.24 ;
      RECT 116.41 222.48 116.76 222.64 ;
      RECT 116.41 225.88 116.76 226.04 ;
      RECT 116.41 229.28 116.76 229.44 ;
      RECT 116.41 232.68 116.76 232.84 ;
      RECT 116.41 236.08 116.76 236.24 ;
      RECT 116.41 239.48 116.76 239.64 ;
      RECT 116.41 242.88 116.76 243.04 ;
      RECT 116.41 246.28 116.76 246.44 ;
      RECT 116.41 249.68 116.76 249.84 ;
      RECT 116.41 253.08 116.76 253.24 ;
      RECT 116.41 256.48 116.76 256.64 ;
      RECT 116.41 259.88 116.76 260.04 ;
      RECT 116.41 263.28 116.76 263.44 ;
      RECT 116.41 266.68 116.76 266.84 ;
      RECT 116.41 270.08 116.76 270.24 ;
      RECT 116.41 273.48 116.76 273.64 ;
      RECT 116.41 276.88 116.76 277.04 ;
      RECT 116.41 280.28 116.76 280.44 ;
      RECT 116.41 283.68 116.76 283.84 ;
      RECT 116.41 287.08 116.76 287.24 ;
      RECT 116.41 290.48 116.76 290.64 ;
      RECT 116.41 293.88 116.76 294.04 ;
      RECT 116.41 297.28 116.76 297.44 ;
      RECT 116.41 300.68 116.76 300.84 ;
      RECT 116.41 304.08 116.76 304.24 ;
      RECT 116.41 307.48 116.76 307.64 ;
      RECT 116.41 310.88 116.76 311.04 ;
      RECT 116.41 314.28 116.76 314.44 ;
      RECT 116.41 317.68 116.76 317.84 ;
      RECT 116.41 321.08 116.76 321.24 ;
      RECT 116.41 324.48 116.76 324.64 ;
      RECT 116.41 327.88 116.76 328.04 ;
      RECT 116.41 331.28 116.76 331.44 ;
      RECT 116.41 334.68 116.76 334.84 ;
      RECT 116.41 338.08 116.76 338.24 ;
      RECT 116.41 341.48 116.76 341.64 ;
      RECT 116.41 344.88 116.76 345.04 ;
      RECT 116.41 348.28 116.76 348.44 ;
      RECT 116.41 351.68 116.76 351.84 ;
      RECT 116.41 355.08 116.76 355.24 ;
      RECT 116.41 358.48 116.76 358.64 ;
      RECT 116.41 361.88 116.76 362.04 ;
      RECT 116.41 365.28 116.76 365.44 ;
      RECT 116.41 368.68 116.76 368.84 ;
      RECT 116.41 372.08 116.76 372.24 ;
      RECT 116.41 375.48 116.76 375.64 ;
      RECT 116.41 378.88 116.76 379.04 ;
      RECT 116.41 382.28 116.76 382.44 ;
      RECT 116.41 385.68 116.76 385.84 ;
      RECT 116.41 389.08 116.76 389.24 ;
      RECT 116.41 392.48 116.76 392.64 ;
      RECT 116.41 395.88 116.76 396.04 ;
      RECT 116.41 399.28 116.76 399.44 ;
      RECT 116.41 402.68 116.76 402.84 ;
      RECT 116.41 406.08 116.76 406.24 ;
      RECT 116.41 409.48 116.76 409.64 ;
      RECT 116.41 412.88 116.76 413.04 ;
      RECT 116.41 416.28 116.76 416.44 ;
      RECT 116.41 419.68 116.76 419.84 ;
      RECT 116.41 423.08 116.76 423.24 ;
      RECT 116.41 426.48 116.76 426.64 ;
      RECT 116.41 429.88 116.76 430.04 ;
      RECT 116.41 433.28 116.76 433.44 ;
      RECT 116.41 436.68 116.76 436.84 ;
      RECT 116.41 440.08 116.76 440.24 ;
      RECT 116.41 443.48 116.76 443.64 ;
      RECT 116.41 446.88 116.76 447.04 ;
      RECT 116.41 450.28 116.76 450.44 ;
      RECT 116.41 453.68 116.76 453.84 ;
      RECT 116.41 457.08 116.76 457.24 ;
      RECT 116.41 460.48 116.76 460.64 ;
      RECT 116.41 463.88 116.76 464.04 ;
      RECT 116.41 467.28 116.76 467.44 ;
      RECT 116.41 470.68 116.76 470.84 ;
      RECT 116.41 474.08 116.76 474.24 ;
      RECT 116.41 477.48 116.76 477.64 ;
      RECT 116.41 480.88 116.76 481.04 ;
      RECT 116.41 484.28 116.76 484.44 ;
      RECT 116.41 487.68 116.76 487.84 ;
      RECT 116.41 491.08 116.76 491.24 ;
      RECT 116.41 494.48 116.76 494.64 ;
      RECT 116.41 497.88 116.76 498.04 ;
      RECT 116.41 9.61 116.57 14.44 ;
      RECT 115.84 76.28 116.25 76.44 ;
      RECT 115.84 83.08 116.25 83.24 ;
      RECT 115.84 89.88 116.25 90.04 ;
      RECT 115.84 96.68 116.25 96.84 ;
      RECT 115.84 103.48 116.25 103.64 ;
      RECT 115.84 110.28 116.25 110.44 ;
      RECT 115.84 117.08 116.25 117.24 ;
      RECT 115.84 123.88 116.25 124.04 ;
      RECT 115.84 130.68 116.25 130.84 ;
      RECT 115.84 137.48 116.25 137.64 ;
      RECT 115.84 144.28 116.25 144.44 ;
      RECT 115.84 151.08 116.25 151.24 ;
      RECT 115.84 157.88 116.25 158.04 ;
      RECT 115.84 164.68 116.25 164.84 ;
      RECT 115.84 171.48 116.25 171.64 ;
      RECT 115.84 178.28 116.25 178.44 ;
      RECT 115.84 185.08 116.25 185.24 ;
      RECT 115.84 191.88 116.25 192.04 ;
      RECT 115.84 198.68 116.25 198.84 ;
      RECT 115.84 205.48 116.25 205.64 ;
      RECT 115.93 12.63 116.09 17.44 ;
      RECT 115.93 17.6 116.09 20.88 ;
      RECT 115.93 32.85 116.09 36.97 ;
      RECT 115.93 40.73 116.09 41.55 ;
      RECT 115.93 60.41 116.09 64 ;
      RECT 115.45 9.61 115.61 14.44 ;
      RECT 115.24 37.58 115.43 38.41 ;
      RECT 115.11 38.57 115.27 40.5 ;
      RECT 114.82 37.58 114.99 38.41 ;
      RECT 114.71 17.46 114.87 20.88 ;
      RECT 114.71 61.17 114.87 64.59 ;
      RECT 113.97 23.99 114.65 24.21 ;
      RECT 113.97 57.84 114.65 58.06 ;
      RECT 114.14 7.04 114.46 7.36 ;
      RECT 111.21 510.54 114.01 510.94 ;
      RECT 113.64 37.58 113.92 38.41 ;
      RECT 113.75 17.46 113.91 20.88 ;
      RECT 113.75 61.17 113.91 64.59 ;
      RECT 111.61 6.24 113.59 6.84 ;
      RECT 113.35 38.57 113.51 40.5 ;
      RECT 113.19 37.58 113.48 38.41 ;
      RECT 113.27 30.54 113.43 32.2 ;
      RECT 113.27 50.09 113.43 51.7 ;
      RECT 113.01 9.61 113.17 14.44 ;
      RECT 112.5 23.97 112.72 24.48 ;
      RECT 112.5 57.58 112.72 58.08 ;
      RECT 112.53 12.63 112.69 17.44 ;
      RECT 112.53 31.09 112.69 36.97 ;
      RECT 112.53 40.73 112.69 41.55 ;
      RECT 112.53 45.65 112.69 51.3 ;
      RECT 111.74 37.58 112.03 38.41 ;
      RECT 111.79 30.54 111.95 32.2 ;
      RECT 111.79 50.09 111.95 51.7 ;
      RECT 111.71 38.57 111.87 40.5 ;
      RECT 111.3 37.58 111.58 38.41 ;
      RECT 111.31 14.52 111.47 16.86 ;
      RECT 111.31 17.46 111.47 20.88 ;
      RECT 111.31 61.17 111.47 64.59 ;
      RECT 110.57 23.99 111.25 24.21 ;
      RECT 110.57 57.84 111.25 58.06 ;
      RECT 110.35 14.52 110.51 16.86 ;
      RECT 110.35 17.46 110.51 20.88 ;
      RECT 110.35 61.17 110.51 64.59 ;
      RECT 110.23 37.58 110.4 38.41 ;
      RECT 108.23 6.24 110.21 6.84 ;
      RECT 109.95 38.57 110.11 40.5 ;
      RECT 109.79 37.58 109.98 38.41 ;
      RECT 109.13 12.63 109.29 17.44 ;
      RECT 109.13 17.6 109.29 20.88 ;
      RECT 109.13 32.85 109.29 36.97 ;
      RECT 109.13 40.73 109.29 41.55 ;
      RECT 109.13 60.41 109.29 64 ;
      RECT 107.81 510.36 108.91 510.94 ;
      RECT 108.65 9.61 108.81 14.44 ;
      RECT 108.44 37.58 108.63 38.41 ;
      RECT 108.31 38.57 108.47 40.5 ;
      RECT 108.02 37.58 108.19 38.41 ;
      RECT 107.91 17.46 108.07 20.88 ;
      RECT 107.91 61.17 108.07 64.59 ;
      RECT 107.8 505.32 107.96 505.88 ;
      RECT 107.17 23.99 107.85 24.21 ;
      RECT 107.17 57.84 107.85 58.06 ;
      RECT 107.34 7.04 107.66 7.36 ;
      RECT 107.02 505.32 107.18 505.88 ;
      RECT 106.84 37.58 107.12 38.41 ;
      RECT 106.95 17.46 107.11 20.88 ;
      RECT 106.95 61.17 107.11 64.59 ;
      RECT 104.83 6.24 106.79 6.84 ;
      RECT 106.55 38.57 106.71 40.5 ;
      RECT 106.39 37.58 106.68 38.41 ;
      RECT 106.47 30.54 106.63 32.2 ;
      RECT 106.47 50.09 106.63 51.7 ;
      RECT 106.21 9.61 106.37 14.44 ;
      RECT 105.7 23.97 105.92 24.48 ;
      RECT 105.7 57.58 105.92 58.08 ;
      RECT 105.73 12.63 105.89 17.44 ;
      RECT 105.73 31.09 105.89 36.97 ;
      RECT 105.73 40.73 105.89 41.55 ;
      RECT 105.73 45.65 105.89 51.3 ;
      RECT 102.71 73.1 105.51 75.96 ;
      RECT 102.71 76.76 105.51 79.62 ;
      RECT 102.71 79.9 105.51 82.76 ;
      RECT 102.71 86.7 105.51 89.56 ;
      RECT 102.71 90.36 105.51 93.22 ;
      RECT 102.71 93.5 105.51 96.36 ;
      RECT 102.71 100.3 105.51 103.16 ;
      RECT 102.71 103.96 105.51 106.82 ;
      RECT 102.71 107.1 105.51 109.96 ;
      RECT 102.71 113.9 105.51 116.76 ;
      RECT 102.71 117.56 105.51 120.42 ;
      RECT 102.71 120.7 105.51 123.56 ;
      RECT 102.71 127.5 105.51 130.36 ;
      RECT 102.71 131.16 105.51 134.02 ;
      RECT 102.71 134.3 105.51 137.16 ;
      RECT 102.71 141.1 105.51 143.96 ;
      RECT 102.71 144.76 105.51 147.62 ;
      RECT 102.71 147.9 105.51 150.76 ;
      RECT 102.71 154.7 105.51 157.56 ;
      RECT 102.71 158.36 105.51 161.22 ;
      RECT 102.71 161.5 105.51 164.36 ;
      RECT 102.71 168.3 105.51 171.16 ;
      RECT 102.71 171.96 105.51 174.82 ;
      RECT 102.71 175.1 105.51 177.96 ;
      RECT 102.71 181.9 105.51 184.76 ;
      RECT 102.71 185.56 105.51 188.42 ;
      RECT 102.71 188.7 105.51 191.56 ;
      RECT 102.71 195.5 105.51 198.36 ;
      RECT 102.71 199.16 105.51 202.02 ;
      RECT 102.71 202.3 105.51 205.16 ;
      RECT 102.71 209.1 105.51 211.96 ;
      RECT 102.71 212.76 105.51 215.62 ;
      RECT 102.71 215.9 105.51 218.76 ;
      RECT 102.71 222.7 105.51 225.56 ;
      RECT 102.71 226.36 105.51 229.22 ;
      RECT 102.71 229.5 105.51 232.36 ;
      RECT 102.71 236.3 105.51 239.16 ;
      RECT 102.71 239.96 105.51 242.82 ;
      RECT 102.71 243.1 105.51 245.96 ;
      RECT 102.71 249.9 105.51 252.76 ;
      RECT 102.71 253.56 105.51 256.42 ;
      RECT 102.71 256.7 105.51 259.56 ;
      RECT 102.71 263.5 105.51 266.36 ;
      RECT 102.71 267.16 105.51 270.02 ;
      RECT 102.71 270.3 105.51 273.16 ;
      RECT 102.71 277.1 105.51 279.96 ;
      RECT 102.71 280.76 105.51 283.62 ;
      RECT 102.71 283.9 105.51 286.76 ;
      RECT 102.71 290.7 105.51 293.56 ;
      RECT 102.71 294.36 105.51 297.22 ;
      RECT 102.71 297.5 105.51 300.36 ;
      RECT 102.71 304.3 105.51 307.16 ;
      RECT 102.71 307.96 105.51 310.82 ;
      RECT 102.71 311.1 105.51 313.96 ;
      RECT 102.71 317.9 105.51 320.76 ;
      RECT 102.71 321.56 105.51 324.42 ;
      RECT 102.71 324.7 105.51 327.56 ;
      RECT 102.71 331.5 105.51 334.36 ;
      RECT 102.71 335.16 105.51 338.02 ;
      RECT 102.71 338.3 105.51 341.16 ;
      RECT 102.71 345.1 105.51 347.96 ;
      RECT 102.71 348.76 105.51 351.62 ;
      RECT 102.71 351.9 105.51 354.76 ;
      RECT 102.71 358.7 105.51 361.56 ;
      RECT 102.71 362.36 105.51 365.22 ;
      RECT 102.71 365.5 105.51 368.36 ;
      RECT 102.71 372.3 105.51 375.16 ;
      RECT 102.71 375.96 105.51 378.82 ;
      RECT 102.71 379.1 105.51 381.96 ;
      RECT 102.71 385.9 105.51 388.76 ;
      RECT 102.71 389.56 105.51 392.42 ;
      RECT 102.71 392.7 105.51 395.56 ;
      RECT 102.71 399.5 105.51 402.36 ;
      RECT 102.71 403.16 105.51 406.02 ;
      RECT 102.71 406.3 105.51 409.16 ;
      RECT 102.71 413.1 105.51 415.96 ;
      RECT 102.71 416.76 105.51 419.62 ;
      RECT 102.71 419.9 105.51 422.76 ;
      RECT 102.71 426.7 105.51 429.56 ;
      RECT 102.71 430.36 105.51 433.22 ;
      RECT 102.71 433.5 105.51 436.36 ;
      RECT 102.71 440.3 105.51 443.16 ;
      RECT 102.71 443.96 105.51 446.82 ;
      RECT 102.71 447.1 105.51 449.96 ;
      RECT 102.71 453.9 105.51 456.76 ;
      RECT 102.71 457.56 105.51 460.42 ;
      RECT 102.71 460.7 105.51 463.56 ;
      RECT 102.71 467.5 105.51 470.36 ;
      RECT 102.71 471.16 105.51 474.02 ;
      RECT 102.71 474.3 105.51 477.16 ;
      RECT 102.71 481.1 105.51 483.96 ;
      RECT 102.71 484.76 105.51 487.62 ;
      RECT 102.71 487.9 105.51 490.76 ;
      RECT 102.71 494.7 105.51 497.56 ;
      RECT 102.71 498.36 105.51 501.22 ;
      RECT 102.71 501.5 105.51 504.36 ;
      RECT 104.41 510.36 105.51 510.94 ;
      RECT 105.25 9.61 105.41 14.44 ;
      RECT 104.94 37.58 105.23 38.41 ;
      RECT 104.99 30.54 105.15 32.2 ;
      RECT 104.99 50.09 105.15 51.7 ;
      RECT 104.91 38.57 105.07 40.5 ;
      RECT 104.5 37.58 104.78 38.41 ;
      RECT 104.51 17.46 104.67 20.88 ;
      RECT 104.51 61.17 104.67 64.59 ;
      RECT 104.4 505.32 104.56 505.88 ;
      RECT 103.77 23.99 104.45 24.21 ;
      RECT 103.77 57.84 104.45 58.06 ;
      RECT 103.96 7.04 104.28 7.36 ;
      RECT 103.62 505.32 103.78 505.88 ;
      RECT 103.55 17.46 103.71 20.88 ;
      RECT 103.55 61.17 103.71 64.59 ;
      RECT 103.43 37.58 103.6 38.41 ;
      RECT 101.43 6.24 103.39 6.84 ;
      RECT 103.15 38.57 103.31 40.5 ;
      RECT 102.99 37.58 103.18 38.41 ;
      RECT 102.81 9.61 102.97 14.44 ;
      RECT 102.33 12.63 102.49 17.44 ;
      RECT 102.33 17.6 102.49 20.88 ;
      RECT 102.33 32.85 102.49 36.97 ;
      RECT 102.33 40.73 102.49 41.55 ;
      RECT 102.33 60.41 102.49 64 ;
      RECT 99.31 73.1 102.11 75.96 ;
      RECT 99.31 76.76 102.11 79.62 ;
      RECT 99.31 79.9 102.11 82.76 ;
      RECT 99.31 86.7 102.11 89.56 ;
      RECT 99.31 90.36 102.11 93.22 ;
      RECT 99.31 93.5 102.11 96.36 ;
      RECT 99.31 100.3 102.11 103.16 ;
      RECT 99.31 103.96 102.11 106.82 ;
      RECT 99.31 107.1 102.11 109.96 ;
      RECT 99.31 113.9 102.11 116.76 ;
      RECT 99.31 117.56 102.11 120.42 ;
      RECT 99.31 120.7 102.11 123.56 ;
      RECT 99.31 127.5 102.11 130.36 ;
      RECT 99.31 131.16 102.11 134.02 ;
      RECT 99.31 134.3 102.11 137.16 ;
      RECT 99.31 141.1 102.11 143.96 ;
      RECT 99.31 144.76 102.11 147.62 ;
      RECT 99.31 147.9 102.11 150.76 ;
      RECT 99.31 154.7 102.11 157.56 ;
      RECT 99.31 158.36 102.11 161.22 ;
      RECT 99.31 161.5 102.11 164.36 ;
      RECT 99.31 168.3 102.11 171.16 ;
      RECT 99.31 171.96 102.11 174.82 ;
      RECT 99.31 175.1 102.11 177.96 ;
      RECT 99.31 181.9 102.11 184.76 ;
      RECT 99.31 185.56 102.11 188.42 ;
      RECT 99.31 188.7 102.11 191.56 ;
      RECT 99.31 195.5 102.11 198.36 ;
      RECT 99.31 199.16 102.11 202.02 ;
      RECT 99.31 202.3 102.11 205.16 ;
      RECT 99.31 209.1 102.11 211.96 ;
      RECT 99.31 212.76 102.11 215.62 ;
      RECT 99.31 215.9 102.11 218.76 ;
      RECT 99.31 222.7 102.11 225.56 ;
      RECT 99.31 226.36 102.11 229.22 ;
      RECT 99.31 229.5 102.11 232.36 ;
      RECT 99.31 236.3 102.11 239.16 ;
      RECT 99.31 239.96 102.11 242.82 ;
      RECT 99.31 243.1 102.11 245.96 ;
      RECT 99.31 249.9 102.11 252.76 ;
      RECT 99.31 253.56 102.11 256.42 ;
      RECT 99.31 256.7 102.11 259.56 ;
      RECT 99.31 263.5 102.11 266.36 ;
      RECT 99.31 267.16 102.11 270.02 ;
      RECT 99.31 270.3 102.11 273.16 ;
      RECT 99.31 277.1 102.11 279.96 ;
      RECT 99.31 280.76 102.11 283.62 ;
      RECT 99.31 283.9 102.11 286.76 ;
      RECT 99.31 290.7 102.11 293.56 ;
      RECT 99.31 294.36 102.11 297.22 ;
      RECT 99.31 297.5 102.11 300.36 ;
      RECT 99.31 304.3 102.11 307.16 ;
      RECT 99.31 307.96 102.11 310.82 ;
      RECT 99.31 311.1 102.11 313.96 ;
      RECT 99.31 317.9 102.11 320.76 ;
      RECT 99.31 321.56 102.11 324.42 ;
      RECT 99.31 324.7 102.11 327.56 ;
      RECT 99.31 331.5 102.11 334.36 ;
      RECT 99.31 335.16 102.11 338.02 ;
      RECT 99.31 338.3 102.11 341.16 ;
      RECT 99.31 345.1 102.11 347.96 ;
      RECT 99.31 348.76 102.11 351.62 ;
      RECT 99.31 351.9 102.11 354.76 ;
      RECT 99.31 358.7 102.11 361.56 ;
      RECT 99.31 362.36 102.11 365.22 ;
      RECT 99.31 365.5 102.11 368.36 ;
      RECT 99.31 372.3 102.11 375.16 ;
      RECT 99.31 375.96 102.11 378.82 ;
      RECT 99.31 379.1 102.11 381.96 ;
      RECT 99.31 385.9 102.11 388.76 ;
      RECT 99.31 389.56 102.11 392.42 ;
      RECT 99.31 392.7 102.11 395.56 ;
      RECT 99.31 399.5 102.11 402.36 ;
      RECT 99.31 403.16 102.11 406.02 ;
      RECT 99.31 406.3 102.11 409.16 ;
      RECT 99.31 413.1 102.11 415.96 ;
      RECT 99.31 416.76 102.11 419.62 ;
      RECT 99.31 419.9 102.11 422.76 ;
      RECT 99.31 426.7 102.11 429.56 ;
      RECT 99.31 430.36 102.11 433.22 ;
      RECT 99.31 433.5 102.11 436.36 ;
      RECT 99.31 440.3 102.11 443.16 ;
      RECT 99.31 443.96 102.11 446.82 ;
      RECT 99.31 447.1 102.11 449.96 ;
      RECT 99.31 453.9 102.11 456.76 ;
      RECT 99.31 457.56 102.11 460.42 ;
      RECT 99.31 460.7 102.11 463.56 ;
      RECT 99.31 467.5 102.11 470.36 ;
      RECT 99.31 471.16 102.11 474.02 ;
      RECT 99.31 474.3 102.11 477.16 ;
      RECT 99.31 481.1 102.11 483.96 ;
      RECT 99.31 484.76 102.11 487.62 ;
      RECT 99.31 487.9 102.11 490.76 ;
      RECT 99.31 494.7 102.11 497.56 ;
      RECT 99.31 498.36 102.11 501.22 ;
      RECT 99.31 501.5 102.11 504.36 ;
      RECT 101.01 510.36 102.11 510.94 ;
      RECT 101.85 9.61 102.01 14.44 ;
      RECT 101.64 37.58 101.83 38.41 ;
      RECT 101.51 38.57 101.67 40.5 ;
      RECT 101.22 37.58 101.39 38.41 ;
      RECT 101.11 17.46 101.27 20.88 ;
      RECT 101.11 61.17 101.27 64.59 ;
      RECT 101 505.32 101.16 505.88 ;
      RECT 100.37 23.99 101.05 24.21 ;
      RECT 100.37 57.84 101.05 58.06 ;
      RECT 100.54 7.04 100.86 7.36 ;
      RECT 100.22 505.32 100.38 505.88 ;
      RECT 100.04 37.58 100.32 38.41 ;
      RECT 100.15 17.46 100.31 20.88 ;
      RECT 100.15 61.17 100.31 64.59 ;
      RECT 98.01 6.24 99.99 6.84 ;
      RECT 99.75 38.57 99.91 40.5 ;
      RECT 99.59 37.58 99.88 38.41 ;
      RECT 99.67 30.54 99.83 32.2 ;
      RECT 99.67 50.09 99.83 51.7 ;
      RECT 99.41 9.61 99.57 14.44 ;
      RECT 98.9 23.97 99.12 24.48 ;
      RECT 98.9 57.58 99.12 58.08 ;
      RECT 98.93 12.63 99.09 17.44 ;
      RECT 98.93 31.09 99.09 36.97 ;
      RECT 98.93 40.73 99.09 41.55 ;
      RECT 98.93 45.65 99.09 51.3 ;
      RECT 95.91 73.1 98.71 75.96 ;
      RECT 95.91 76.76 98.71 79.62 ;
      RECT 95.91 79.9 98.71 82.76 ;
      RECT 95.91 86.7 98.71 89.56 ;
      RECT 95.91 90.36 98.71 93.22 ;
      RECT 95.91 93.5 98.71 96.36 ;
      RECT 95.91 100.3 98.71 103.16 ;
      RECT 95.91 103.96 98.71 106.82 ;
      RECT 95.91 107.1 98.71 109.96 ;
      RECT 95.91 113.9 98.71 116.76 ;
      RECT 95.91 117.56 98.71 120.42 ;
      RECT 95.91 120.7 98.71 123.56 ;
      RECT 95.91 127.5 98.71 130.36 ;
      RECT 95.91 131.16 98.71 134.02 ;
      RECT 95.91 134.3 98.71 137.16 ;
      RECT 95.91 141.1 98.71 143.96 ;
      RECT 95.91 144.76 98.71 147.62 ;
      RECT 95.91 147.9 98.71 150.76 ;
      RECT 95.91 154.7 98.71 157.56 ;
      RECT 95.91 158.36 98.71 161.22 ;
      RECT 95.91 161.5 98.71 164.36 ;
      RECT 95.91 168.3 98.71 171.16 ;
      RECT 95.91 171.96 98.71 174.82 ;
      RECT 95.91 175.1 98.71 177.96 ;
      RECT 95.91 181.9 98.71 184.76 ;
      RECT 95.91 185.56 98.71 188.42 ;
      RECT 95.91 188.7 98.71 191.56 ;
      RECT 95.91 195.5 98.71 198.36 ;
      RECT 95.91 199.16 98.71 202.02 ;
      RECT 95.91 202.3 98.71 205.16 ;
      RECT 95.91 209.1 98.71 211.96 ;
      RECT 95.91 212.76 98.71 215.62 ;
      RECT 95.91 215.9 98.71 218.76 ;
      RECT 95.91 222.7 98.71 225.56 ;
      RECT 95.91 226.36 98.71 229.22 ;
      RECT 95.91 229.5 98.71 232.36 ;
      RECT 95.91 236.3 98.71 239.16 ;
      RECT 95.91 239.96 98.71 242.82 ;
      RECT 95.91 243.1 98.71 245.96 ;
      RECT 95.91 249.9 98.71 252.76 ;
      RECT 95.91 253.56 98.71 256.42 ;
      RECT 95.91 256.7 98.71 259.56 ;
      RECT 95.91 263.5 98.71 266.36 ;
      RECT 95.91 267.16 98.71 270.02 ;
      RECT 95.91 270.3 98.71 273.16 ;
      RECT 95.91 277.1 98.71 279.96 ;
      RECT 95.91 280.76 98.71 283.62 ;
      RECT 95.91 283.9 98.71 286.76 ;
      RECT 95.91 290.7 98.71 293.56 ;
      RECT 95.91 294.36 98.71 297.22 ;
      RECT 95.91 297.5 98.71 300.36 ;
      RECT 95.91 304.3 98.71 307.16 ;
      RECT 95.91 307.96 98.71 310.82 ;
      RECT 95.91 311.1 98.71 313.96 ;
      RECT 95.91 317.9 98.71 320.76 ;
      RECT 95.91 321.56 98.71 324.42 ;
      RECT 95.91 324.7 98.71 327.56 ;
      RECT 95.91 331.5 98.71 334.36 ;
      RECT 95.91 335.16 98.71 338.02 ;
      RECT 95.91 338.3 98.71 341.16 ;
      RECT 95.91 345.1 98.71 347.96 ;
      RECT 95.91 348.76 98.71 351.62 ;
      RECT 95.91 351.9 98.71 354.76 ;
      RECT 95.91 358.7 98.71 361.56 ;
      RECT 95.91 362.36 98.71 365.22 ;
      RECT 95.91 365.5 98.71 368.36 ;
      RECT 95.91 372.3 98.71 375.16 ;
      RECT 95.91 375.96 98.71 378.82 ;
      RECT 95.91 379.1 98.71 381.96 ;
      RECT 95.91 385.9 98.71 388.76 ;
      RECT 95.91 389.56 98.71 392.42 ;
      RECT 95.91 392.7 98.71 395.56 ;
      RECT 95.91 399.5 98.71 402.36 ;
      RECT 95.91 403.16 98.71 406.02 ;
      RECT 95.91 406.3 98.71 409.16 ;
      RECT 95.91 413.1 98.71 415.96 ;
      RECT 95.91 416.76 98.71 419.62 ;
      RECT 95.91 419.9 98.71 422.76 ;
      RECT 95.91 426.7 98.71 429.56 ;
      RECT 95.91 430.36 98.71 433.22 ;
      RECT 95.91 433.5 98.71 436.36 ;
      RECT 95.91 440.3 98.71 443.16 ;
      RECT 95.91 443.96 98.71 446.82 ;
      RECT 95.91 447.1 98.71 449.96 ;
      RECT 95.91 453.9 98.71 456.76 ;
      RECT 95.91 457.56 98.71 460.42 ;
      RECT 95.91 460.7 98.71 463.56 ;
      RECT 95.91 467.5 98.71 470.36 ;
      RECT 95.91 471.16 98.71 474.02 ;
      RECT 95.91 474.3 98.71 477.16 ;
      RECT 95.91 481.1 98.71 483.96 ;
      RECT 95.91 484.76 98.71 487.62 ;
      RECT 95.91 487.9 98.71 490.76 ;
      RECT 95.91 494.7 98.71 497.56 ;
      RECT 95.91 498.36 98.71 501.22 ;
      RECT 95.91 501.5 98.71 504.36 ;
      RECT 97.61 510.36 98.71 510.94 ;
      RECT 98.14 37.58 98.43 38.41 ;
      RECT 98.19 30.54 98.35 32.2 ;
      RECT 98.19 50.09 98.35 51.7 ;
      RECT 98.11 38.57 98.27 40.5 ;
      RECT 97.7 37.58 97.98 38.41 ;
      RECT 97.71 14.52 97.87 16.86 ;
      RECT 97.71 17.46 97.87 20.88 ;
      RECT 97.71 61.17 97.87 64.59 ;
      RECT 97.6 505.32 97.76 505.88 ;
      RECT 96.97 23.99 97.65 24.21 ;
      RECT 96.97 57.84 97.65 58.06 ;
      RECT 96.82 505.32 96.98 505.88 ;
      RECT 96.75 14.52 96.91 16.86 ;
      RECT 96.75 17.46 96.91 20.88 ;
      RECT 96.75 61.17 96.91 64.59 ;
      RECT 96.63 37.58 96.8 38.41 ;
      RECT 94.63 6.24 96.61 6.84 ;
      RECT 96.35 38.57 96.51 40.5 ;
      RECT 96.19 37.58 96.38 38.41 ;
      RECT 95.53 12.63 95.69 17.44 ;
      RECT 95.53 17.6 95.69 20.88 ;
      RECT 95.53 32.85 95.69 36.97 ;
      RECT 95.53 40.73 95.69 41.55 ;
      RECT 95.53 60.41 95.69 64 ;
      RECT 92.51 69.86 95.31 72.66 ;
      RECT 92.51 73.1 95.31 75.96 ;
      RECT 92.51 76.76 95.31 79.62 ;
      RECT 92.51 79.9 95.31 82.76 ;
      RECT 92.51 83.56 95.31 86.42 ;
      RECT 92.51 86.7 95.31 89.56 ;
      RECT 92.51 90.36 95.31 93.22 ;
      RECT 92.51 93.5 95.31 96.36 ;
      RECT 92.51 97.16 95.31 100.02 ;
      RECT 92.51 100.3 95.31 103.16 ;
      RECT 92.51 103.96 95.31 106.82 ;
      RECT 92.51 107.1 95.31 109.96 ;
      RECT 92.51 110.76 95.31 113.62 ;
      RECT 92.51 113.9 95.31 116.76 ;
      RECT 92.51 117.56 95.31 120.42 ;
      RECT 92.51 120.7 95.31 123.56 ;
      RECT 92.51 124.36 95.31 127.22 ;
      RECT 92.51 127.5 95.31 130.36 ;
      RECT 92.51 131.16 95.31 134.02 ;
      RECT 92.51 134.3 95.31 137.16 ;
      RECT 92.51 137.96 95.31 140.82 ;
      RECT 92.51 141.1 95.31 143.96 ;
      RECT 92.51 144.76 95.31 147.62 ;
      RECT 92.51 147.9 95.31 150.76 ;
      RECT 92.51 151.56 95.31 154.42 ;
      RECT 92.51 154.7 95.31 157.56 ;
      RECT 92.51 158.36 95.31 161.22 ;
      RECT 92.51 161.5 95.31 164.36 ;
      RECT 92.51 165.16 95.31 168.02 ;
      RECT 92.51 168.3 95.31 171.16 ;
      RECT 92.51 171.96 95.31 174.82 ;
      RECT 92.51 175.1 95.31 177.96 ;
      RECT 92.51 178.66 95.31 181.46 ;
      RECT 92.51 181.9 95.31 184.76 ;
      RECT 92.51 185.56 95.31 188.42 ;
      RECT 92.51 188.7 95.31 191.56 ;
      RECT 92.51 192.36 95.31 195.22 ;
      RECT 92.51 195.5 95.31 198.36 ;
      RECT 92.51 199.16 95.31 202.02 ;
      RECT 92.51 202.3 95.31 205.16 ;
      RECT 92.51 205.96 95.31 208.82 ;
      RECT 92.51 209.1 95.31 211.96 ;
      RECT 92.51 212.76 95.31 215.62 ;
      RECT 92.51 215.9 95.31 218.76 ;
      RECT 92.51 219.56 95.31 222.42 ;
      RECT 92.51 222.7 95.31 225.56 ;
      RECT 92.51 226.36 95.31 229.22 ;
      RECT 92.51 229.5 95.31 232.36 ;
      RECT 92.51 233.16 95.31 236.02 ;
      RECT 92.51 236.3 95.31 239.16 ;
      RECT 92.51 239.96 95.31 242.82 ;
      RECT 92.51 243.1 95.31 245.96 ;
      RECT 92.51 246.76 95.31 249.62 ;
      RECT 92.51 249.9 95.31 252.76 ;
      RECT 92.51 253.56 95.31 256.42 ;
      RECT 92.51 256.7 95.31 259.56 ;
      RECT 92.51 260.36 95.31 263.22 ;
      RECT 92.51 263.5 95.31 266.36 ;
      RECT 92.51 267.16 95.31 270.02 ;
      RECT 92.51 270.3 95.31 273.16 ;
      RECT 92.51 273.96 95.31 276.82 ;
      RECT 92.51 277.1 95.31 279.96 ;
      RECT 92.51 280.76 95.31 283.62 ;
      RECT 92.51 283.9 95.31 286.76 ;
      RECT 92.51 287.46 95.31 290.26 ;
      RECT 92.51 290.7 95.31 293.56 ;
      RECT 92.51 294.36 95.31 297.22 ;
      RECT 92.51 297.5 95.31 300.36 ;
      RECT 92.51 301.16 95.31 304.02 ;
      RECT 92.51 304.3 95.31 307.16 ;
      RECT 92.51 307.96 95.31 310.82 ;
      RECT 92.51 311.1 95.31 313.96 ;
      RECT 92.51 314.76 95.31 317.62 ;
      RECT 92.51 317.9 95.31 320.76 ;
      RECT 92.51 321.56 95.31 324.42 ;
      RECT 92.51 324.7 95.31 327.56 ;
      RECT 92.51 328.36 95.31 331.22 ;
      RECT 92.51 331.5 95.31 334.36 ;
      RECT 92.51 335.16 95.31 338.02 ;
      RECT 92.51 338.3 95.31 341.16 ;
      RECT 92.51 341.96 95.31 344.82 ;
      RECT 92.51 345.1 95.31 347.96 ;
      RECT 92.51 348.76 95.31 351.62 ;
      RECT 92.51 351.9 95.31 354.76 ;
      RECT 92.51 355.56 95.31 358.42 ;
      RECT 92.51 358.7 95.31 361.56 ;
      RECT 92.51 362.36 95.31 365.22 ;
      RECT 92.51 365.5 95.31 368.36 ;
      RECT 92.51 369.16 95.31 372.02 ;
      RECT 92.51 372.3 95.31 375.16 ;
      RECT 92.51 375.96 95.31 378.82 ;
      RECT 92.51 379.1 95.31 381.96 ;
      RECT 92.51 382.76 95.31 385.62 ;
      RECT 92.51 385.9 95.31 388.76 ;
      RECT 92.51 389.56 95.31 392.42 ;
      RECT 92.51 392.7 95.31 395.56 ;
      RECT 92.51 396.26 95.31 399.06 ;
      RECT 92.51 399.5 95.31 402.36 ;
      RECT 92.51 403.16 95.31 406.02 ;
      RECT 92.51 406.3 95.31 409.16 ;
      RECT 92.51 409.96 95.31 412.82 ;
      RECT 92.51 413.1 95.31 415.96 ;
      RECT 92.51 416.76 95.31 419.62 ;
      RECT 92.51 419.9 95.31 422.76 ;
      RECT 92.51 423.56 95.31 426.42 ;
      RECT 92.51 426.7 95.31 429.56 ;
      RECT 92.51 430.36 95.31 433.22 ;
      RECT 92.51 433.5 95.31 436.36 ;
      RECT 92.51 437.16 95.31 440.02 ;
      RECT 92.51 440.3 95.31 443.16 ;
      RECT 92.51 443.96 95.31 446.82 ;
      RECT 92.51 447.1 95.31 449.96 ;
      RECT 92.51 450.76 95.31 453.62 ;
      RECT 92.51 453.9 95.31 456.76 ;
      RECT 92.51 457.56 95.31 460.42 ;
      RECT 92.51 460.7 95.31 463.56 ;
      RECT 92.51 464.36 95.31 467.22 ;
      RECT 92.51 467.5 95.31 470.36 ;
      RECT 92.51 471.16 95.31 474.02 ;
      RECT 92.51 474.3 95.31 477.16 ;
      RECT 92.51 477.96 95.31 480.82 ;
      RECT 92.51 481.1 95.31 483.96 ;
      RECT 92.51 484.76 95.31 487.62 ;
      RECT 92.51 487.9 95.31 490.76 ;
      RECT 92.51 491.56 95.31 494.42 ;
      RECT 92.51 494.7 95.31 497.56 ;
      RECT 92.51 498.36 95.31 501.22 ;
      RECT 92.51 501.5 95.31 504.36 ;
      RECT 94.21 510.36 95.31 510.94 ;
      RECT 95.05 9.61 95.21 14.44 ;
      RECT 94.84 37.58 95.03 38.41 ;
      RECT 94.71 38.57 94.87 40.5 ;
      RECT 94.42 37.58 94.59 38.41 ;
      RECT 94.31 17.46 94.47 20.88 ;
      RECT 94.31 61.17 94.47 64.59 ;
      RECT 94.2 505.32 94.36 505.88 ;
      RECT 93.57 23.99 94.25 24.21 ;
      RECT 93.57 57.84 94.25 58.06 ;
      RECT 93.74 7.04 94.06 7.36 ;
      RECT 93.42 505.32 93.58 505.88 ;
      RECT 93.24 37.58 93.52 38.41 ;
      RECT 93.35 17.46 93.51 20.88 ;
      RECT 93.35 61.17 93.51 64.59 ;
      RECT 91.23 6.24 93.19 6.84 ;
      RECT 92.95 38.57 93.11 40.5 ;
      RECT 92.79 37.58 93.08 38.41 ;
      RECT 92.87 30.54 93.03 32.2 ;
      RECT 92.87 50.09 93.03 51.7 ;
      RECT 92.61 9.61 92.77 14.44 ;
      RECT 92.1 23.97 92.32 24.48 ;
      RECT 92.1 57.58 92.32 58.08 ;
      RECT 92.13 12.63 92.29 17.44 ;
      RECT 92.13 31.09 92.29 36.97 ;
      RECT 92.13 40.73 92.29 41.55 ;
      RECT 92.13 45.65 92.29 51.3 ;
      RECT 89.11 69.85 91.91 72.65 ;
      RECT 89.11 73.1 91.91 75.96 ;
      RECT 89.11 76.76 91.91 79.62 ;
      RECT 89.11 79.9 91.91 82.76 ;
      RECT 89.11 83.56 91.91 86.42 ;
      RECT 89.11 86.7 91.91 89.56 ;
      RECT 89.11 90.36 91.91 93.22 ;
      RECT 89.11 93.5 91.91 96.36 ;
      RECT 89.11 97.16 91.91 100.02 ;
      RECT 89.11 100.3 91.91 103.16 ;
      RECT 89.11 103.96 91.91 106.82 ;
      RECT 89.11 107.1 91.91 109.96 ;
      RECT 89.11 110.76 91.91 113.62 ;
      RECT 89.11 113.9 91.91 116.76 ;
      RECT 89.11 117.56 91.91 120.42 ;
      RECT 89.11 120.7 91.91 123.56 ;
      RECT 89.11 124.36 91.91 127.22 ;
      RECT 89.11 127.5 91.91 130.36 ;
      RECT 89.11 131.16 91.91 134.02 ;
      RECT 89.11 134.3 91.91 137.16 ;
      RECT 89.11 137.96 91.91 140.82 ;
      RECT 89.11 141.1 91.91 143.96 ;
      RECT 89.11 144.76 91.91 147.62 ;
      RECT 89.11 147.9 91.91 150.76 ;
      RECT 89.11 151.56 91.91 154.42 ;
      RECT 89.11 154.7 91.91 157.56 ;
      RECT 89.11 158.36 91.91 161.22 ;
      RECT 89.11 161.5 91.91 164.36 ;
      RECT 89.11 165.16 91.91 168.02 ;
      RECT 89.11 168.3 91.91 171.16 ;
      RECT 89.11 171.96 91.91 174.82 ;
      RECT 89.11 175.1 91.91 177.96 ;
      RECT 89.11 178.65 91.91 181.45 ;
      RECT 89.11 181.9 91.91 184.76 ;
      RECT 89.11 185.56 91.91 188.42 ;
      RECT 89.11 188.7 91.91 191.56 ;
      RECT 89.11 192.36 91.91 195.22 ;
      RECT 89.11 195.5 91.91 198.36 ;
      RECT 89.11 199.16 91.91 202.02 ;
      RECT 89.11 202.3 91.91 205.16 ;
      RECT 89.11 205.96 91.91 208.82 ;
      RECT 89.11 209.1 91.91 211.96 ;
      RECT 89.11 212.76 91.91 215.62 ;
      RECT 89.11 215.9 91.91 218.76 ;
      RECT 89.11 219.56 91.91 222.42 ;
      RECT 89.11 222.7 91.91 225.56 ;
      RECT 89.11 226.36 91.91 229.22 ;
      RECT 89.11 229.5 91.91 232.36 ;
      RECT 89.11 233.16 91.91 236.02 ;
      RECT 89.11 236.3 91.91 239.16 ;
      RECT 89.11 239.96 91.91 242.82 ;
      RECT 89.11 243.1 91.91 245.96 ;
      RECT 89.11 246.76 91.91 249.62 ;
      RECT 89.11 249.9 91.91 252.76 ;
      RECT 89.11 253.56 91.91 256.42 ;
      RECT 89.11 256.7 91.91 259.56 ;
      RECT 89.11 260.36 91.91 263.22 ;
      RECT 89.11 263.5 91.91 266.36 ;
      RECT 89.11 267.16 91.91 270.02 ;
      RECT 89.11 270.3 91.91 273.16 ;
      RECT 89.11 273.96 91.91 276.82 ;
      RECT 89.11 277.1 91.91 279.96 ;
      RECT 89.11 280.76 91.91 283.62 ;
      RECT 89.11 283.9 91.91 286.76 ;
      RECT 89.11 287.45 91.91 290.25 ;
      RECT 89.11 290.7 91.91 293.56 ;
      RECT 89.11 294.36 91.91 297.22 ;
      RECT 89.11 297.5 91.91 300.36 ;
      RECT 89.11 301.16 91.91 304.02 ;
      RECT 89.11 304.3 91.91 307.16 ;
      RECT 89.11 307.96 91.91 310.82 ;
      RECT 89.11 311.1 91.91 313.96 ;
      RECT 89.11 314.76 91.91 317.62 ;
      RECT 89.11 317.9 91.91 320.76 ;
      RECT 89.11 321.56 91.91 324.42 ;
      RECT 89.11 324.7 91.91 327.56 ;
      RECT 89.11 328.36 91.91 331.22 ;
      RECT 89.11 331.5 91.91 334.36 ;
      RECT 89.11 335.16 91.91 338.02 ;
      RECT 89.11 338.3 91.91 341.16 ;
      RECT 89.11 341.96 91.91 344.82 ;
      RECT 89.11 345.1 91.91 347.96 ;
      RECT 89.11 348.76 91.91 351.62 ;
      RECT 89.11 351.9 91.91 354.76 ;
      RECT 89.11 355.56 91.91 358.42 ;
      RECT 89.11 358.7 91.91 361.56 ;
      RECT 89.11 362.36 91.91 365.22 ;
      RECT 89.11 365.5 91.91 368.36 ;
      RECT 89.11 369.16 91.91 372.02 ;
      RECT 89.11 372.3 91.91 375.16 ;
      RECT 89.11 375.96 91.91 378.82 ;
      RECT 89.11 379.1 91.91 381.96 ;
      RECT 89.11 382.76 91.91 385.62 ;
      RECT 89.11 385.9 91.91 388.76 ;
      RECT 89.11 389.56 91.91 392.42 ;
      RECT 89.11 392.7 91.91 395.56 ;
      RECT 89.11 396.25 91.91 399.05 ;
      RECT 89.11 399.5 91.91 402.36 ;
      RECT 89.11 403.16 91.91 406.02 ;
      RECT 89.11 406.3 91.91 409.16 ;
      RECT 89.11 409.96 91.91 412.82 ;
      RECT 89.11 413.1 91.91 415.96 ;
      RECT 89.11 416.76 91.91 419.62 ;
      RECT 89.11 419.9 91.91 422.76 ;
      RECT 89.11 423.56 91.91 426.42 ;
      RECT 89.11 426.7 91.91 429.56 ;
      RECT 89.11 430.36 91.91 433.22 ;
      RECT 89.11 433.5 91.91 436.36 ;
      RECT 89.11 437.16 91.91 440.02 ;
      RECT 89.11 440.3 91.91 443.16 ;
      RECT 89.11 443.96 91.91 446.82 ;
      RECT 89.11 447.1 91.91 449.96 ;
      RECT 89.11 450.76 91.91 453.62 ;
      RECT 89.11 453.9 91.91 456.76 ;
      RECT 89.11 457.56 91.91 460.42 ;
      RECT 89.11 460.7 91.91 463.56 ;
      RECT 89.11 464.36 91.91 467.22 ;
      RECT 89.11 467.5 91.91 470.36 ;
      RECT 89.11 471.16 91.91 474.02 ;
      RECT 89.11 474.3 91.91 477.16 ;
      RECT 89.11 477.96 91.91 480.82 ;
      RECT 89.11 481.1 91.91 483.96 ;
      RECT 89.11 484.76 91.91 487.62 ;
      RECT 89.11 487.9 91.91 490.76 ;
      RECT 89.11 491.56 91.91 494.42 ;
      RECT 89.11 494.7 91.91 497.56 ;
      RECT 89.11 498.36 91.91 501.22 ;
      RECT 89.11 501.5 91.91 504.36 ;
      RECT 90.81 510.36 91.91 510.94 ;
      RECT 91.65 9.61 91.81 14.44 ;
      RECT 91.34 37.58 91.63 38.41 ;
      RECT 91.39 30.54 91.55 32.2 ;
      RECT 91.39 50.09 91.55 51.7 ;
      RECT 91.31 38.57 91.47 40.5 ;
      RECT 90.9 37.58 91.18 38.41 ;
      RECT 90.91 17.46 91.07 20.88 ;
      RECT 90.91 61.17 91.07 64.59 ;
      RECT 90.8 505.32 90.96 505.88 ;
      RECT 90.17 23.99 90.85 24.21 ;
      RECT 90.17 57.84 90.85 58.06 ;
      RECT 90.36 7.04 90.68 7.36 ;
      RECT 90.02 505.32 90.18 505.88 ;
      RECT 89.95 17.46 90.11 20.88 ;
      RECT 89.95 61.17 90.11 64.59 ;
      RECT 89.83 37.58 90 38.41 ;
      RECT 88.81 6.24 89.79 6.84 ;
      RECT 89.55 38.57 89.71 40.5 ;
      RECT 89.39 37.58 89.58 38.41 ;
      RECT 89.21 9.61 89.37 14.44 ;
      RECT 88.73 12.63 88.89 17.44 ;
      RECT 88.73 17.6 88.89 20.88 ;
      RECT 88.73 32.85 88.89 36.97 ;
      RECT 88.73 40.73 88.89 41.55 ;
      RECT 88.73 60.41 88.89 64 ;
      RECT 87.81 510.36 88.61 510.94 ;
      RECT 87.21 6.24 88.01 6.64 ;
      RECT 85.41 6.24 86.71 6.84 ;
      RECT 86.31 36.22 86.51 36.95 ;
      RECT 86.33 29.32 86.49 34.08 ;
      RECT 86.33 39.34 86.49 46.59 ;
      RECT 86.33 47.59 86.49 51.92 ;
      RECT 86.33 52.64 86.49 56.5 ;
      RECT 86.01 47.88 86.17 51.16 ;
      RECT 85.85 57.79 86.01 62.72 ;
      RECT 85.61 29.97 85.77 32.28 ;
      RECT 85.61 35.23 85.77 36.31 ;
      RECT 85.61 37.11 85.77 38.19 ;
      RECT 85.61 41.14 85.77 43.45 ;
      RECT 77.69 15.46 85.53 16.9 ;
      RECT 85.37 57.79 85.53 62.72 ;
      RECT 85.01 56.99 85.41 57.29 ;
      RECT 85.13 29.97 85.29 34.08 ;
      RECT 85.13 39.34 85.29 43.45 ;
      RECT 85.05 48.24 85.21 50.5 ;
      RECT 84.89 57.79 85.05 67.9 ;
      RECT 83.03 6.24 85.01 6.84 ;
      RECT 83.01 510.54 85.01 510.94 ;
      RECT 84.65 29.97 84.81 32.28 ;
      RECT 84.65 35.23 84.81 36.31 ;
      RECT 84.65 37.11 84.81 38.19 ;
      RECT 84.65 41.14 84.81 43.45 ;
      RECT 78.59 21.67 84.63 21.95 ;
      RECT 83.91 36.21 84.11 36.95 ;
      RECT 83.93 29.32 84.09 34.08 ;
      RECT 83.93 39.34 84.09 46.59 ;
      RECT 83.93 47.59 84.09 51.11 ;
      RECT 83.93 51.34 84.09 53.67 ;
      RECT 83.93 54.16 84.09 56.5 ;
      RECT 83.21 29.97 83.37 32.28 ;
      RECT 83.21 35.23 83.37 36.31 ;
      RECT 83.21 37.11 83.37 38.19 ;
      RECT 83.21 41.14 83.37 43.45 ;
      RECT 82.97 57.79 83.13 67.9 ;
      RECT 82.61 56.99 83.01 57.29 ;
      RECT 82.81 48.24 82.97 50.5 ;
      RECT 82.73 29.97 82.89 34.08 ;
      RECT 82.73 39.34 82.89 43.45 ;
      RECT 82.49 57.79 82.65 62.72 ;
      RECT 80.63 6.24 82.61 6.84 ;
      RECT 82.25 29.97 82.41 32.28 ;
      RECT 82.25 35.23 82.41 36.31 ;
      RECT 82.25 37.11 82.41 38.19 ;
      RECT 82.25 41.14 82.41 43.45 ;
      RECT 82.01 57.79 82.17 62.72 ;
      RECT 81.85 47.88 82.01 51.16 ;
      RECT 81.33 9.36 81.89 9.52 ;
      RECT 81.33 11.3 81.89 11.46 ;
      RECT 81.33 14.68 81.89 14.84 ;
      RECT 81.33 19.63 81.89 19.79 ;
      RECT 81.51 36.21 81.71 36.95 ;
      RECT 81.53 29.32 81.69 34.08 ;
      RECT 81.53 39.34 81.69 46.59 ;
      RECT 81.53 47.59 81.69 51.92 ;
      RECT 81.53 52.64 81.69 56.5 ;
      RECT 81.21 47.88 81.37 51.16 ;
      RECT 81.05 57.79 81.21 62.72 ;
      RECT 80.81 29.97 80.97 32.28 ;
      RECT 80.81 35.23 80.97 36.31 ;
      RECT 80.81 37.11 80.97 38.19 ;
      RECT 80.81 41.14 80.97 43.45 ;
      RECT 80.57 57.79 80.73 62.72 ;
      RECT 80.21 56.99 80.61 57.29 ;
      RECT 80.33 29.97 80.49 34.08 ;
      RECT 80.33 39.34 80.49 43.45 ;
      RECT 80.25 48.24 80.41 50.5 ;
      RECT 80.09 57.79 80.25 67.9 ;
      RECT 78.23 6.24 80.21 6.84 ;
      RECT 78.21 510.54 80.21 510.94 ;
      RECT 79.85 29.97 80.01 32.28 ;
      RECT 79.85 35.23 80.01 36.31 ;
      RECT 79.85 37.11 80.01 38.19 ;
      RECT 79.85 41.14 80.01 43.45 ;
      RECT 79.11 36.21 79.31 36.95 ;
      RECT 79.13 29.32 79.29 34.08 ;
      RECT 79.13 39.34 79.29 46.59 ;
      RECT 79.13 47.59 79.29 51.11 ;
      RECT 79.13 51.34 79.29 53.67 ;
      RECT 79.13 54.16 79.29 56.5 ;
      RECT 78.41 29.97 78.57 32.28 ;
      RECT 78.41 35.23 78.57 36.31 ;
      RECT 78.41 37.11 78.57 38.19 ;
      RECT 78.41 41.14 78.57 43.45 ;
      RECT 78.17 57.79 78.33 67.9 ;
      RECT 77.81 56.99 78.21 57.29 ;
      RECT 78.01 48.24 78.17 50.5 ;
      RECT 77.93 29.97 78.09 34.08 ;
      RECT 77.93 39.34 78.09 43.45 ;
      RECT 77.69 57.79 77.85 62.72 ;
      RECT 75.81 6.24 77.81 6.84 ;
      RECT 77.45 29.97 77.61 32.28 ;
      RECT 77.45 35.23 77.61 36.31 ;
      RECT 77.45 37.11 77.61 38.19 ;
      RECT 77.45 41.14 77.61 43.45 ;
      RECT 77.21 57.79 77.37 62.72 ;
      RECT 77.05 47.88 77.21 51.16 ;
      RECT 76.71 36.21 76.91 36.95 ;
      RECT 76.73 21.45 76.89 24.52 ;
      RECT 76.73 29.32 76.89 34.08 ;
      RECT 76.73 39.34 76.89 46.59 ;
      RECT 76.73 47.59 76.89 51.92 ;
      RECT 76.73 52.64 76.89 56.5 ;
      RECT 76.06 8.96 76.57 9.17 ;
      RECT 76.41 47.83 76.57 51.16 ;
      RECT 76.27 15.09 76.55 15.41 ;
      RECT 76.25 57.79 76.41 62.72 ;
      RECT 76.05 12.28 76.37 12.76 ;
      RECT 76.09 21.73 76.25 22.33 ;
      RECT 76.09 22.49 76.25 23.06 ;
      RECT 76.01 29.97 76.17 32.28 ;
      RECT 76.01 35.23 76.17 36.31 ;
      RECT 76.01 37.11 76.17 38.19 ;
      RECT 76.01 41.14 76.17 43.45 ;
      RECT 75.77 57.79 75.93 62.72 ;
      RECT 75.41 56.99 75.81 57.29 ;
      RECT 74.63 13.4 75.75 13.56 ;
      RECT 75.53 29.97 75.69 34.08 ;
      RECT 75.53 39.34 75.69 43.45 ;
      RECT 75.52 26.68 75.68 28.17 ;
      RECT 75.45 48.24 75.61 50.5 ;
      RECT 75.25 10.76 75.57 11.16 ;
      RECT 74.83 10 75.55 10.18 ;
      RECT 75.29 57.79 75.45 67.9 ;
      RECT 73.44 6.24 75.41 6.84 ;
      RECT 73.41 510.54 75.41 510.94 ;
      RECT 75.05 29.97 75.21 32.28 ;
      RECT 75.05 35.23 75.21 36.31 ;
      RECT 75.05 37.11 75.21 38.19 ;
      RECT 75.05 41.14 75.21 43.45 ;
      RECT 74.74 17 74.9 18.12 ;
      RECT 74.31 36.21 74.51 36.95 ;
      RECT 74.33 29.32 74.49 34.08 ;
      RECT 74.33 39.34 74.49 46.59 ;
      RECT 74.33 47.59 74.49 51.11 ;
      RECT 74.33 51.34 74.49 53.67 ;
      RECT 74.33 54.16 74.49 56.5 ;
      RECT 74.01 23.54 74.45 23.81 ;
      RECT 74.1 15.33 74.26 15.89 ;
      RECT 73.54 28.33 74.1 28.49 ;
      RECT 73.61 25.51 73.85 26.2 ;
      RECT 73.61 29.97 73.77 32.28 ;
      RECT 73.61 35.23 73.77 36.31 ;
      RECT 73.61 37.11 73.77 38.19 ;
      RECT 73.61 41.14 73.77 43.45 ;
      RECT 73.37 57.79 73.53 67.9 ;
      RECT 73.01 56.99 73.41 57.29 ;
      RECT 73.22 16.21 73.38 18.62 ;
      RECT 73.21 48.24 73.37 50.5 ;
      RECT 73.13 29.97 73.29 34.08 ;
      RECT 73.13 39.34 73.29 43.45 ;
      RECT 73.07 14.84 73.23 16.05 ;
      RECT 72.89 57.79 73.05 62.72 ;
      RECT 71.51 6.24 73.01 6.84 ;
      RECT 72.65 29.97 72.81 32.28 ;
      RECT 72.65 35.23 72.81 36.31 ;
      RECT 72.65 37.11 72.81 38.19 ;
      RECT 72.65 41.14 72.81 43.45 ;
      RECT 72.41 57.79 72.57 62.72 ;
      RECT 72.19 19.63 72.51 20.04 ;
      RECT 72.25 47.88 72.41 51.16 ;
      RECT 71.75 13.8 72.31 13.96 ;
      RECT 71.63 13.32 72.11 13.56 ;
      RECT 71.91 36.21 72.11 36.95 ;
      RECT 71.93 26.38 72.09 27.85 ;
      RECT 71.93 29.32 72.09 34.08 ;
      RECT 71.93 39.34 72.09 46.59 ;
      RECT 71.93 47.59 72.09 51.92 ;
      RECT 71.93 52.64 72.09 56.5 ;
      RECT 71.61 47.88 71.77 51.16 ;
      RECT 71.21 16.47 71.63 17.1 ;
      RECT 71.45 57.79 71.61 62.72 ;
      RECT 71.21 29.97 71.37 32.28 ;
      RECT 71.21 35.23 71.37 36.31 ;
      RECT 71.21 37.11 71.37 38.19 ;
      RECT 71.21 41.14 71.37 43.45 ;
      RECT 70.97 57.79 71.13 62.72 ;
      RECT 70.61 56.99 71.01 57.29 ;
      RECT 70.73 29.97 70.89 34.08 ;
      RECT 70.73 39.34 70.89 43.45 ;
      RECT 70.65 48.24 70.81 50.5 ;
      RECT 70.49 57.79 70.65 67.9 ;
      RECT 68.61 510.54 70.61 510.94 ;
      RECT 69.92 28.33 70.48 28.49 ;
      RECT 70.17 25.51 70.41 26.2 ;
      RECT 70.25 29.97 70.41 32.28 ;
      RECT 70.25 35.23 70.41 36.31 ;
      RECT 70.25 37.11 70.41 38.19 ;
      RECT 70.25 41.14 70.41 43.45 ;
      RECT 69.11 6.24 70.11 6.84 ;
      RECT 69.57 23.54 70.01 23.81 ;
      RECT 69.51 36.21 69.71 36.95 ;
      RECT 69.53 29.32 69.69 34.08 ;
      RECT 69.53 39.34 69.69 46.59 ;
      RECT 69.53 47.59 69.69 51.11 ;
      RECT 69.53 51.34 69.69 53.67 ;
      RECT 69.53 54.16 69.69 56.5 ;
      RECT 69.33 21.85 69.49 22.91 ;
      RECT 69.3 7.58 69.46 8.64 ;
      RECT 69.26 20.65 69.42 21.69 ;
      RECT 67.95 16.8 68.97 17.08 ;
      RECT 68.81 29.97 68.97 32.28 ;
      RECT 68.81 35.23 68.97 36.31 ;
      RECT 68.81 37.11 68.97 38.19 ;
      RECT 68.81 41.14 68.97 43.45 ;
      RECT 68.49 15.32 68.89 15.64 ;
      RECT 68.57 57.79 68.73 67.9 ;
      RECT 68.21 56.99 68.61 57.29 ;
      RECT 68.42 8.04 68.58 8.6 ;
      RECT 68.41 48.24 68.57 50.5 ;
      RECT 67.95 16.12 68.51 16.28 ;
      RECT 68.34 26.68 68.5 28.17 ;
      RECT 68.33 29.97 68.49 34.08 ;
      RECT 68.33 39.34 68.49 43.45 ;
      RECT 68.09 11.52 68.25 13.07 ;
      RECT 68.09 57.79 68.25 62.72 ;
      RECT 67.85 29.97 68.01 32.28 ;
      RECT 67.85 35.23 68.01 36.31 ;
      RECT 67.85 37.11 68.01 38.19 ;
      RECT 67.85 41.14 68.01 43.45 ;
      RECT 67.73 13.11 67.89 13.67 ;
      RECT 67.61 57.79 67.77 62.72 ;
      RECT 66.81 6.24 67.61 6.84 ;
      RECT 67.45 47.88 67.61 51.16 ;
      RECT 67.11 36.21 67.31 36.95 ;
      RECT 67.13 21.45 67.29 24.52 ;
      RECT 67.13 29.32 67.29 34.08 ;
      RECT 67.13 39.34 67.29 46.59 ;
      RECT 67.13 47.59 67.29 51.92 ;
      RECT 67.13 52.64 67.29 56.5 ;
      RECT 66.81 47.88 66.97 51.16 ;
      RECT 66.65 57.79 66.81 62.72 ;
      RECT 66.53 13.11 66.69 13.67 ;
      RECT 66.41 29.97 66.57 32.28 ;
      RECT 66.41 35.23 66.57 36.31 ;
      RECT 66.41 37.11 66.57 38.19 ;
      RECT 66.41 41.14 66.57 43.45 ;
      RECT 65.91 16.12 66.47 16.28 ;
      RECT 65.45 16.8 66.47 17.08 ;
      RECT 66.17 11.52 66.33 13.07 ;
      RECT 66.17 57.79 66.33 62.72 ;
      RECT 65.81 56.99 66.21 57.29 ;
      RECT 65.93 29.97 66.09 34.08 ;
      RECT 65.93 39.34 66.09 43.45 ;
      RECT 65.92 26.68 66.08 28.17 ;
      RECT 65.85 48.24 66.01 50.5 ;
      RECT 65.84 8.04 66 8.6 ;
      RECT 65.53 15.32 65.93 15.64 ;
      RECT 65.69 57.79 65.85 67.9 ;
      RECT 63.81 510.54 65.81 510.94 ;
      RECT 65.45 29.97 65.61 32.28 ;
      RECT 65.45 35.23 65.61 36.31 ;
      RECT 65.45 37.11 65.61 38.19 ;
      RECT 65.45 41.14 65.61 43.45 ;
      RECT 64.31 6.24 65.31 6.84 ;
      RECT 65 20.65 65.16 21.69 ;
      RECT 64.96 7.58 65.12 8.64 ;
      RECT 64.93 21.85 65.09 22.91 ;
      RECT 64.71 36.21 64.91 36.95 ;
      RECT 64.73 29.32 64.89 34.08 ;
      RECT 64.73 39.34 64.89 46.59 ;
      RECT 64.73 47.59 64.89 51.11 ;
      RECT 64.73 51.34 64.89 53.67 ;
      RECT 64.73 54.16 64.89 56.5 ;
      RECT 64.41 23.54 64.85 23.81 ;
      RECT 63.94 28.33 64.5 28.49 ;
      RECT 64.01 25.51 64.25 26.2 ;
      RECT 64.01 29.97 64.17 32.28 ;
      RECT 64.01 35.23 64.17 36.31 ;
      RECT 64.01 37.11 64.17 38.19 ;
      RECT 64.01 41.14 64.17 43.45 ;
      RECT 63.77 57.79 63.93 67.9 ;
      RECT 63.41 56.99 63.81 57.29 ;
      RECT 63.61 48.24 63.77 50.5 ;
      RECT 63.53 29.97 63.69 34.08 ;
      RECT 63.53 39.34 63.69 43.45 ;
      RECT 63.29 57.79 63.45 62.72 ;
      RECT 62.79 16.47 63.21 17.1 ;
      RECT 63.05 29.97 63.21 32.28 ;
      RECT 63.05 35.23 63.21 36.31 ;
      RECT 63.05 37.11 63.21 38.19 ;
      RECT 63.05 41.14 63.21 43.45 ;
      RECT 62.81 57.79 62.97 62.72 ;
      RECT 61.41 6.24 62.91 6.84 ;
      RECT 62.65 47.88 62.81 51.16 ;
      RECT 62.31 13.32 62.79 13.56 ;
      RECT 62.11 13.8 62.67 13.96 ;
      RECT 62.31 36.21 62.51 36.95 ;
      RECT 62.33 26.38 62.49 27.85 ;
      RECT 62.33 29.32 62.49 34.08 ;
      RECT 62.33 39.34 62.49 46.59 ;
      RECT 62.33 47.59 62.49 51.92 ;
      RECT 62.33 52.64 62.49 56.5 ;
      RECT 61.91 19.63 62.23 20.04 ;
      RECT 62.01 47.88 62.17 51.16 ;
      RECT 61.85 57.79 62.01 62.72 ;
      RECT 61.61 29.97 61.77 32.28 ;
      RECT 61.61 35.23 61.77 36.31 ;
      RECT 61.61 37.11 61.77 38.19 ;
      RECT 61.61 41.14 61.77 43.45 ;
      RECT 61.37 57.79 61.53 62.72 ;
      RECT 61.01 56.99 61.41 57.29 ;
      RECT 61.19 14.84 61.35 16.05 ;
      RECT 61.13 29.97 61.29 34.08 ;
      RECT 61.13 39.34 61.29 43.45 ;
      RECT 61.05 48.24 61.21 50.5 ;
      RECT 61.04 16.21 61.2 18.62 ;
      RECT 60.89 57.79 61.05 67.9 ;
      RECT 59.01 510.54 61.01 510.94 ;
      RECT 59.01 6.24 60.98 6.84 ;
      RECT 60.32 28.33 60.88 28.49 ;
      RECT 60.57 25.51 60.81 26.2 ;
      RECT 60.65 29.97 60.81 32.28 ;
      RECT 60.65 35.23 60.81 36.31 ;
      RECT 60.65 37.11 60.81 38.19 ;
      RECT 60.65 41.14 60.81 43.45 ;
      RECT 59.97 23.54 60.41 23.81 ;
      RECT 60.16 15.33 60.32 15.89 ;
      RECT 59.91 36.21 60.11 36.95 ;
      RECT 59.93 29.32 60.09 34.08 ;
      RECT 59.93 39.34 60.09 46.59 ;
      RECT 59.93 47.59 60.09 51.11 ;
      RECT 59.93 51.34 60.09 53.67 ;
      RECT 59.93 54.16 60.09 56.5 ;
      RECT 58.67 13.4 59.79 13.56 ;
      RECT 59.52 17 59.68 18.12 ;
      RECT 58.87 10 59.59 10.18 ;
      RECT 59.21 29.97 59.37 32.28 ;
      RECT 59.21 35.23 59.37 36.31 ;
      RECT 59.21 37.11 59.37 38.19 ;
      RECT 59.21 41.14 59.37 43.45 ;
      RECT 58.85 10.76 59.17 11.16 ;
      RECT 58.97 57.79 59.13 67.9 ;
      RECT 58.61 56.99 59.01 57.29 ;
      RECT 58.81 48.24 58.97 50.5 ;
      RECT 58.74 26.68 58.9 28.17 ;
      RECT 58.73 29.97 58.89 34.08 ;
      RECT 58.73 39.34 58.89 43.45 ;
      RECT 58.49 57.79 58.65 62.72 ;
      RECT 56.61 6.24 58.61 6.84 ;
      RECT 58.25 29.97 58.41 32.28 ;
      RECT 58.25 35.23 58.41 36.31 ;
      RECT 58.25 37.11 58.41 38.19 ;
      RECT 58.25 41.14 58.41 43.45 ;
      RECT 58.05 12.28 58.37 12.76 ;
      RECT 57.85 8.96 58.36 9.17 ;
      RECT 58.17 21.73 58.33 22.33 ;
      RECT 58.17 22.49 58.33 23.06 ;
      RECT 58.01 57.79 58.17 62.72 ;
      RECT 57.87 15.09 58.15 15.41 ;
      RECT 57.85 47.88 58.01 51.16 ;
      RECT 57.51 36.21 57.71 36.95 ;
      RECT 57.53 21.45 57.69 24.52 ;
      RECT 57.53 29.32 57.69 34.08 ;
      RECT 57.53 39.34 57.69 46.59 ;
      RECT 57.53 47.59 57.69 51.92 ;
      RECT 57.53 52.64 57.69 56.5 ;
      RECT 57.21 47.83 57.37 51.16 ;
      RECT 57.05 57.79 57.21 62.72 ;
      RECT 56.81 29.97 56.97 32.28 ;
      RECT 56.81 35.23 56.97 36.31 ;
      RECT 56.81 37.11 56.97 38.19 ;
      RECT 56.81 41.14 56.97 43.45 ;
      RECT 48.89 15.46 56.73 16.9 ;
      RECT 56.57 57.79 56.73 62.72 ;
      RECT 56.21 56.99 56.61 57.29 ;
      RECT 56.33 29.97 56.49 34.08 ;
      RECT 56.33 39.34 56.49 43.45 ;
      RECT 56.25 48.24 56.41 50.5 ;
      RECT 56.09 57.79 56.25 67.9 ;
      RECT 54.21 510.54 56.21 510.94 ;
      RECT 54.21 6.24 56.19 6.84 ;
      RECT 55.85 29.97 56.01 32.28 ;
      RECT 55.85 35.23 56.01 36.31 ;
      RECT 55.85 37.11 56.01 38.19 ;
      RECT 55.85 41.14 56.01 43.45 ;
      RECT 49.79 21.67 55.83 21.95 ;
      RECT 55.11 36.21 55.31 36.95 ;
      RECT 55.13 29.32 55.29 34.08 ;
      RECT 55.13 39.34 55.29 46.59 ;
      RECT 55.13 47.59 55.29 51.11 ;
      RECT 55.13 51.34 55.29 53.67 ;
      RECT 55.13 54.16 55.29 56.5 ;
      RECT 54.41 29.97 54.57 32.28 ;
      RECT 54.41 35.23 54.57 36.31 ;
      RECT 54.41 37.11 54.57 38.19 ;
      RECT 54.41 41.14 54.57 43.45 ;
      RECT 54.17 57.79 54.33 67.9 ;
      RECT 53.81 56.99 54.21 57.29 ;
      RECT 54.01 48.24 54.17 50.5 ;
      RECT 53.93 29.97 54.09 34.08 ;
      RECT 53.93 39.34 54.09 43.45 ;
      RECT 53.69 57.79 53.85 62.72 ;
      RECT 51.81 6.24 53.79 6.84 ;
      RECT 53.45 29.97 53.61 32.28 ;
      RECT 53.45 35.23 53.61 36.31 ;
      RECT 53.45 37.11 53.61 38.19 ;
      RECT 53.45 41.14 53.61 43.45 ;
      RECT 53.21 57.79 53.37 62.72 ;
      RECT 53.05 47.88 53.21 51.16 ;
      RECT 52.53 9.36 53.09 9.52 ;
      RECT 52.53 11.3 53.09 11.46 ;
      RECT 52.53 14.68 53.09 14.84 ;
      RECT 52.53 19.63 53.09 19.79 ;
      RECT 52.71 36.21 52.91 36.95 ;
      RECT 52.73 29.32 52.89 34.08 ;
      RECT 52.73 39.34 52.89 46.59 ;
      RECT 52.73 47.59 52.89 51.92 ;
      RECT 52.73 52.64 52.89 56.5 ;
      RECT 52.41 47.88 52.57 51.16 ;
      RECT 52.25 57.79 52.41 62.72 ;
      RECT 52.01 29.97 52.17 32.28 ;
      RECT 52.01 35.23 52.17 36.31 ;
      RECT 52.01 37.11 52.17 38.19 ;
      RECT 52.01 41.14 52.17 43.45 ;
      RECT 51.77 57.79 51.93 62.72 ;
      RECT 51.41 56.99 51.81 57.29 ;
      RECT 51.53 29.97 51.69 34.08 ;
      RECT 51.53 39.34 51.69 43.45 ;
      RECT 51.45 48.24 51.61 50.5 ;
      RECT 51.29 57.79 51.45 67.9 ;
      RECT 49.41 510.54 51.41 510.94 ;
      RECT 49.41 6.24 51.39 6.84 ;
      RECT 51.05 29.97 51.21 32.28 ;
      RECT 51.05 35.23 51.21 36.31 ;
      RECT 51.05 37.11 51.21 38.19 ;
      RECT 51.05 41.14 51.21 43.45 ;
      RECT 50.31 36.21 50.51 36.95 ;
      RECT 50.33 29.32 50.49 34.08 ;
      RECT 50.33 39.34 50.49 46.59 ;
      RECT 50.33 47.59 50.49 51.11 ;
      RECT 50.33 51.34 50.49 53.67 ;
      RECT 50.33 54.16 50.49 56.5 ;
      RECT 49.61 29.97 49.77 32.28 ;
      RECT 49.61 35.23 49.77 36.31 ;
      RECT 49.61 37.11 49.77 38.19 ;
      RECT 49.61 41.14 49.77 43.45 ;
      RECT 49.37 57.79 49.53 67.9 ;
      RECT 49.01 56.99 49.41 57.29 ;
      RECT 49.21 48.24 49.37 50.5 ;
      RECT 49.13 29.97 49.29 34.08 ;
      RECT 49.13 39.34 49.29 43.45 ;
      RECT 48.89 57.79 49.05 62.72 ;
      RECT 48.65 29.97 48.81 32.28 ;
      RECT 48.65 35.23 48.81 36.31 ;
      RECT 48.65 37.11 48.81 38.19 ;
      RECT 48.65 41.14 48.81 43.45 ;
      RECT 48.41 57.79 48.57 62.72 ;
      RECT 48.25 47.88 48.41 51.16 ;
      RECT 47.91 36.21 48.11 36.95 ;
      RECT 47.93 29.32 48.09 34.08 ;
      RECT 47.93 39.34 48.09 46.59 ;
      RECT 47.93 47.59 48.09 51.92 ;
      RECT 47.93 52.64 48.09 56.5 ;
      RECT 47.31 36.11 47.51 58.16 ;
      RECT 47.33 8.48 47.49 10.44 ;
      RECT 47.33 17.36 47.49 17.92 ;
      RECT 47.33 20.74 47.49 27.31 ;
      RECT 46.71 36.22 46.91 36.95 ;
      RECT 46.73 29.32 46.89 34.08 ;
      RECT 46.73 39.34 46.89 46.59 ;
      RECT 46.73 47.59 46.89 51.92 ;
      RECT 46.73 52.64 46.89 56.5 ;
      RECT 46.41 47.88 46.57 51.16 ;
      RECT 46.25 57.79 46.41 62.72 ;
      RECT 46.01 29.97 46.17 32.28 ;
      RECT 46.01 35.23 46.17 36.31 ;
      RECT 46.01 37.11 46.17 38.19 ;
      RECT 46.01 41.14 46.17 43.45 ;
      RECT 38.09 15.46 45.93 16.9 ;
      RECT 45.77 57.79 45.93 62.72 ;
      RECT 45.41 56.99 45.81 57.29 ;
      RECT 45.53 29.97 45.69 34.08 ;
      RECT 45.53 39.34 45.69 43.45 ;
      RECT 45.45 48.24 45.61 50.5 ;
      RECT 45.29 57.79 45.45 67.9 ;
      RECT 43.43 6.24 45.41 6.84 ;
      RECT 43.41 510.54 45.41 510.94 ;
      RECT 45.05 29.97 45.21 32.28 ;
      RECT 45.05 35.23 45.21 36.31 ;
      RECT 45.05 37.11 45.21 38.19 ;
      RECT 45.05 41.14 45.21 43.45 ;
      RECT 38.99 21.67 45.03 21.95 ;
      RECT 44.31 36.21 44.51 36.95 ;
      RECT 44.33 29.32 44.49 34.08 ;
      RECT 44.33 39.34 44.49 46.59 ;
      RECT 44.33 47.59 44.49 51.11 ;
      RECT 44.33 51.34 44.49 53.67 ;
      RECT 44.33 54.16 44.49 56.5 ;
      RECT 43.61 29.97 43.77 32.28 ;
      RECT 43.61 35.23 43.77 36.31 ;
      RECT 43.61 37.11 43.77 38.19 ;
      RECT 43.61 41.14 43.77 43.45 ;
      RECT 43.37 57.79 43.53 67.9 ;
      RECT 43.01 56.99 43.41 57.29 ;
      RECT 43.21 48.24 43.37 50.5 ;
      RECT 43.13 29.97 43.29 34.08 ;
      RECT 43.13 39.34 43.29 43.45 ;
      RECT 42.89 57.79 43.05 62.72 ;
      RECT 41.03 6.24 43.01 6.84 ;
      RECT 42.65 29.97 42.81 32.28 ;
      RECT 42.65 35.23 42.81 36.31 ;
      RECT 42.65 37.11 42.81 38.19 ;
      RECT 42.65 41.14 42.81 43.45 ;
      RECT 42.41 57.79 42.57 62.72 ;
      RECT 42.25 47.88 42.41 51.16 ;
      RECT 41.73 9.36 42.29 9.52 ;
      RECT 41.73 11.3 42.29 11.46 ;
      RECT 41.73 14.68 42.29 14.84 ;
      RECT 41.73 19.63 42.29 19.79 ;
      RECT 41.91 36.21 42.11 36.95 ;
      RECT 41.93 29.32 42.09 34.08 ;
      RECT 41.93 39.34 42.09 46.59 ;
      RECT 41.93 47.59 42.09 51.92 ;
      RECT 41.93 52.64 42.09 56.5 ;
      RECT 41.61 47.88 41.77 51.16 ;
      RECT 41.45 57.79 41.61 62.72 ;
      RECT 41.21 29.97 41.37 32.28 ;
      RECT 41.21 35.23 41.37 36.31 ;
      RECT 41.21 37.11 41.37 38.19 ;
      RECT 41.21 41.14 41.37 43.45 ;
      RECT 40.97 57.79 41.13 62.72 ;
      RECT 40.61 56.99 41.01 57.29 ;
      RECT 40.73 29.97 40.89 34.08 ;
      RECT 40.73 39.34 40.89 43.45 ;
      RECT 40.65 48.24 40.81 50.5 ;
      RECT 40.49 57.79 40.65 67.9 ;
      RECT 38.63 6.24 40.61 6.84 ;
      RECT 38.61 510.54 40.61 510.94 ;
      RECT 40.25 29.97 40.41 32.28 ;
      RECT 40.25 35.23 40.41 36.31 ;
      RECT 40.25 37.11 40.41 38.19 ;
      RECT 40.25 41.14 40.41 43.45 ;
      RECT 39.51 36.21 39.71 36.95 ;
      RECT 39.53 29.32 39.69 34.08 ;
      RECT 39.53 39.34 39.69 46.59 ;
      RECT 39.53 47.59 39.69 51.11 ;
      RECT 39.53 51.34 39.69 53.67 ;
      RECT 39.53 54.16 39.69 56.5 ;
      RECT 38.81 29.97 38.97 32.28 ;
      RECT 38.81 35.23 38.97 36.31 ;
      RECT 38.81 37.11 38.97 38.19 ;
      RECT 38.81 41.14 38.97 43.45 ;
      RECT 38.57 57.79 38.73 67.9 ;
      RECT 38.21 56.99 38.61 57.29 ;
      RECT 38.41 48.24 38.57 50.5 ;
      RECT 38.33 29.97 38.49 34.08 ;
      RECT 38.33 39.34 38.49 43.45 ;
      RECT 38.09 57.79 38.25 62.72 ;
      RECT 36.21 6.24 38.21 6.84 ;
      RECT 37.85 29.97 38.01 32.28 ;
      RECT 37.85 35.23 38.01 36.31 ;
      RECT 37.85 37.11 38.01 38.19 ;
      RECT 37.85 41.14 38.01 43.45 ;
      RECT 37.61 57.79 37.77 62.72 ;
      RECT 37.45 47.88 37.61 51.16 ;
      RECT 37.11 36.21 37.31 36.95 ;
      RECT 37.13 21.45 37.29 24.52 ;
      RECT 37.13 29.32 37.29 34.08 ;
      RECT 37.13 39.34 37.29 46.59 ;
      RECT 37.13 47.59 37.29 51.92 ;
      RECT 37.13 52.64 37.29 56.5 ;
      RECT 36.46 8.96 36.97 9.17 ;
      RECT 36.81 47.83 36.97 51.16 ;
      RECT 36.67 15.09 36.95 15.41 ;
      RECT 36.65 57.79 36.81 62.72 ;
      RECT 36.45 12.28 36.77 12.76 ;
      RECT 36.49 21.73 36.65 22.33 ;
      RECT 36.49 22.49 36.65 23.06 ;
      RECT 36.41 29.97 36.57 32.28 ;
      RECT 36.41 35.23 36.57 36.31 ;
      RECT 36.41 37.11 36.57 38.19 ;
      RECT 36.41 41.14 36.57 43.45 ;
      RECT 36.17 57.79 36.33 62.72 ;
      RECT 35.81 56.99 36.21 57.29 ;
      RECT 35.03 13.4 36.15 13.56 ;
      RECT 35.93 29.97 36.09 34.08 ;
      RECT 35.93 39.34 36.09 43.45 ;
      RECT 35.92 26.68 36.08 28.17 ;
      RECT 35.85 48.24 36.01 50.5 ;
      RECT 35.65 10.76 35.97 11.16 ;
      RECT 35.23 10 35.95 10.18 ;
      RECT 35.69 57.79 35.85 67.9 ;
      RECT 33.84 6.24 35.81 6.84 ;
      RECT 33.81 510.54 35.81 510.94 ;
      RECT 35.45 29.97 35.61 32.28 ;
      RECT 35.45 35.23 35.61 36.31 ;
      RECT 35.45 37.11 35.61 38.19 ;
      RECT 35.45 41.14 35.61 43.45 ;
      RECT 35.14 17 35.3 18.12 ;
      RECT 34.71 36.21 34.91 36.95 ;
      RECT 34.73 29.32 34.89 34.08 ;
      RECT 34.73 39.34 34.89 46.59 ;
      RECT 34.73 47.59 34.89 51.11 ;
      RECT 34.73 51.34 34.89 53.67 ;
      RECT 34.73 54.16 34.89 56.5 ;
      RECT 34.41 23.54 34.85 23.81 ;
      RECT 34.5 15.33 34.66 15.89 ;
      RECT 33.94 28.33 34.5 28.49 ;
      RECT 34.01 25.51 34.25 26.2 ;
      RECT 34.01 29.97 34.17 32.28 ;
      RECT 34.01 35.23 34.17 36.31 ;
      RECT 34.01 37.11 34.17 38.19 ;
      RECT 34.01 41.14 34.17 43.45 ;
      RECT 33.77 57.79 33.93 67.9 ;
      RECT 33.41 56.99 33.81 57.29 ;
      RECT 33.62 16.21 33.78 18.62 ;
      RECT 33.61 48.24 33.77 50.5 ;
      RECT 33.53 29.97 33.69 34.08 ;
      RECT 33.53 39.34 33.69 43.45 ;
      RECT 33.47 14.84 33.63 16.05 ;
      RECT 33.29 57.79 33.45 62.72 ;
      RECT 31.91 6.24 33.41 6.84 ;
      RECT 33.05 29.97 33.21 32.28 ;
      RECT 33.05 35.23 33.21 36.31 ;
      RECT 33.05 37.11 33.21 38.19 ;
      RECT 33.05 41.14 33.21 43.45 ;
      RECT 32.81 57.79 32.97 62.72 ;
      RECT 32.59 19.63 32.91 20.04 ;
      RECT 32.65 47.88 32.81 51.16 ;
      RECT 32.15 13.8 32.71 13.96 ;
      RECT 32.03 13.32 32.51 13.56 ;
      RECT 32.31 36.21 32.51 36.95 ;
      RECT 32.33 26.38 32.49 27.85 ;
      RECT 32.33 29.32 32.49 34.08 ;
      RECT 32.33 39.34 32.49 46.59 ;
      RECT 32.33 47.59 32.49 51.92 ;
      RECT 32.33 52.64 32.49 56.5 ;
      RECT 32.01 47.88 32.17 51.16 ;
      RECT 31.61 16.47 32.03 17.1 ;
      RECT 31.85 57.79 32.01 62.72 ;
      RECT 31.61 29.97 31.77 32.28 ;
      RECT 31.61 35.23 31.77 36.31 ;
      RECT 31.61 37.11 31.77 38.19 ;
      RECT 31.61 41.14 31.77 43.45 ;
      RECT 31.37 57.79 31.53 62.72 ;
      RECT 31.01 56.99 31.41 57.29 ;
      RECT 31.13 29.97 31.29 34.08 ;
      RECT 31.13 39.34 31.29 43.45 ;
      RECT 31.05 48.24 31.21 50.5 ;
      RECT 30.89 57.79 31.05 67.9 ;
      RECT 29.01 510.54 31.01 510.94 ;
      RECT 30.32 28.33 30.88 28.49 ;
      RECT 30.57 25.51 30.81 26.2 ;
      RECT 30.65 29.97 30.81 32.28 ;
      RECT 30.65 35.23 30.81 36.31 ;
      RECT 30.65 37.11 30.81 38.19 ;
      RECT 30.65 41.14 30.81 43.45 ;
      RECT 29.51 6.24 30.51 6.84 ;
      RECT 29.97 23.54 30.41 23.81 ;
      RECT 29.91 36.21 30.11 36.95 ;
      RECT 29.93 29.32 30.09 34.08 ;
      RECT 29.93 39.34 30.09 46.59 ;
      RECT 29.93 47.59 30.09 51.11 ;
      RECT 29.93 51.34 30.09 53.67 ;
      RECT 29.93 54.16 30.09 56.5 ;
      RECT 29.73 21.85 29.89 22.91 ;
      RECT 29.7 7.58 29.86 8.64 ;
      RECT 29.66 20.65 29.82 21.69 ;
      RECT 28.35 16.8 29.37 17.08 ;
      RECT 29.21 29.97 29.37 32.28 ;
      RECT 29.21 35.23 29.37 36.31 ;
      RECT 29.21 37.11 29.37 38.19 ;
      RECT 29.21 41.14 29.37 43.45 ;
      RECT 28.89 15.32 29.29 15.64 ;
      RECT 28.97 57.79 29.13 67.9 ;
      RECT 28.61 56.99 29.01 57.29 ;
      RECT 28.82 8.04 28.98 8.6 ;
      RECT 28.81 48.24 28.97 50.5 ;
      RECT 28.35 16.12 28.91 16.28 ;
      RECT 28.74 26.68 28.9 28.17 ;
      RECT 28.73 29.97 28.89 34.08 ;
      RECT 28.73 39.34 28.89 43.45 ;
      RECT 28.49 11.52 28.65 13.07 ;
      RECT 28.49 57.79 28.65 62.72 ;
      RECT 28.25 29.97 28.41 32.28 ;
      RECT 28.25 35.23 28.41 36.31 ;
      RECT 28.25 37.11 28.41 38.19 ;
      RECT 28.25 41.14 28.41 43.45 ;
      RECT 28.13 13.11 28.29 13.67 ;
      RECT 28.01 57.79 28.17 62.72 ;
      RECT 27.21 6.24 28.01 6.84 ;
      RECT 27.85 47.88 28.01 51.16 ;
      RECT 27.51 36.21 27.71 36.95 ;
      RECT 27.53 21.45 27.69 24.52 ;
      RECT 27.53 29.32 27.69 34.08 ;
      RECT 27.53 39.34 27.69 46.59 ;
      RECT 27.53 47.59 27.69 51.92 ;
      RECT 27.53 52.64 27.69 56.5 ;
      RECT 27.21 47.88 27.37 51.16 ;
      RECT 27.05 57.79 27.21 62.72 ;
      RECT 26.93 13.11 27.09 13.67 ;
      RECT 26.81 29.97 26.97 32.28 ;
      RECT 26.81 35.23 26.97 36.31 ;
      RECT 26.81 37.11 26.97 38.19 ;
      RECT 26.81 41.14 26.97 43.45 ;
      RECT 26.31 16.12 26.87 16.28 ;
      RECT 25.85 16.8 26.87 17.08 ;
      RECT 26.57 11.52 26.73 13.07 ;
      RECT 26.57 57.79 26.73 62.72 ;
      RECT 26.21 56.99 26.61 57.29 ;
      RECT 26.33 29.97 26.49 34.08 ;
      RECT 26.33 39.34 26.49 43.45 ;
      RECT 26.32 26.68 26.48 28.17 ;
      RECT 26.25 48.24 26.41 50.5 ;
      RECT 26.24 8.04 26.4 8.6 ;
      RECT 25.93 15.32 26.33 15.64 ;
      RECT 26.09 57.79 26.25 67.9 ;
      RECT 24.21 510.54 26.21 510.94 ;
      RECT 25.85 29.97 26.01 32.28 ;
      RECT 25.85 35.23 26.01 36.31 ;
      RECT 25.85 37.11 26.01 38.19 ;
      RECT 25.85 41.14 26.01 43.45 ;
      RECT 24.71 6.24 25.71 6.84 ;
      RECT 25.4 20.65 25.56 21.69 ;
      RECT 25.36 7.58 25.52 8.64 ;
      RECT 25.33 21.85 25.49 22.91 ;
      RECT 25.11 36.21 25.31 36.95 ;
      RECT 25.13 29.32 25.29 34.08 ;
      RECT 25.13 39.34 25.29 46.59 ;
      RECT 25.13 47.59 25.29 51.11 ;
      RECT 25.13 51.34 25.29 53.67 ;
      RECT 25.13 54.16 25.29 56.5 ;
      RECT 24.81 23.54 25.25 23.81 ;
      RECT 24.34 28.33 24.9 28.49 ;
      RECT 24.41 25.51 24.65 26.2 ;
      RECT 24.41 29.97 24.57 32.28 ;
      RECT 24.41 35.23 24.57 36.31 ;
      RECT 24.41 37.11 24.57 38.19 ;
      RECT 24.41 41.14 24.57 43.45 ;
      RECT 24.17 57.79 24.33 67.9 ;
      RECT 23.81 56.99 24.21 57.29 ;
      RECT 24.01 48.24 24.17 50.5 ;
      RECT 23.93 29.97 24.09 34.08 ;
      RECT 23.93 39.34 24.09 43.45 ;
      RECT 23.69 57.79 23.85 62.72 ;
      RECT 23.19 16.47 23.61 17.1 ;
      RECT 23.45 29.97 23.61 32.28 ;
      RECT 23.45 35.23 23.61 36.31 ;
      RECT 23.45 37.11 23.61 38.19 ;
      RECT 23.45 41.14 23.61 43.45 ;
      RECT 23.21 57.79 23.37 62.72 ;
      RECT 21.81 6.24 23.31 6.84 ;
      RECT 23.05 47.88 23.21 51.16 ;
      RECT 22.71 13.32 23.19 13.56 ;
      RECT 22.51 13.8 23.07 13.96 ;
      RECT 22.71 36.21 22.91 36.95 ;
      RECT 22.73 26.38 22.89 27.85 ;
      RECT 22.73 29.32 22.89 34.08 ;
      RECT 22.73 39.34 22.89 46.59 ;
      RECT 22.73 47.59 22.89 51.92 ;
      RECT 22.73 52.64 22.89 56.5 ;
      RECT 22.31 19.63 22.63 20.04 ;
      RECT 22.41 47.88 22.57 51.16 ;
      RECT 22.25 57.79 22.41 62.72 ;
      RECT 22.01 29.97 22.17 32.28 ;
      RECT 22.01 35.23 22.17 36.31 ;
      RECT 22.01 37.11 22.17 38.19 ;
      RECT 22.01 41.14 22.17 43.45 ;
      RECT 21.77 57.79 21.93 62.72 ;
      RECT 21.41 56.99 21.81 57.29 ;
      RECT 21.59 14.84 21.75 16.05 ;
      RECT 21.53 29.97 21.69 34.08 ;
      RECT 21.53 39.34 21.69 43.45 ;
      RECT 21.45 48.24 21.61 50.5 ;
      RECT 21.44 16.21 21.6 18.62 ;
      RECT 21.29 57.79 21.45 67.9 ;
      RECT 19.81 6.24 21.41 6.84 ;
      RECT 19.41 510.54 21.41 510.94 ;
      RECT 20.72 28.33 21.28 28.49 ;
      RECT 20.97 25.51 21.21 26.2 ;
      RECT 21.05 29.97 21.21 32.28 ;
      RECT 21.05 35.23 21.21 36.31 ;
      RECT 21.05 37.11 21.21 38.19 ;
      RECT 21.05 41.14 21.21 43.45 ;
      RECT 20.37 23.54 20.81 23.81 ;
      RECT 20.56 15.33 20.72 15.89 ;
      RECT 20.31 36.21 20.51 36.95 ;
      RECT 20.33 29.32 20.49 34.08 ;
      RECT 20.33 39.34 20.49 46.59 ;
      RECT 20.33 47.59 20.49 51.11 ;
      RECT 20.33 51.34 20.49 53.67 ;
      RECT 20.33 54.16 20.49 56.5 ;
      RECT 19.07 13.4 20.19 13.56 ;
      RECT 19.92 17 20.08 18.12 ;
      RECT 19.27 10 19.99 10.18 ;
      RECT 19.61 29.97 19.77 32.28 ;
      RECT 19.61 35.23 19.77 36.31 ;
      RECT 19.61 37.11 19.77 38.19 ;
      RECT 19.61 41.14 19.77 43.45 ;
      RECT 19.25 10.76 19.57 11.16 ;
      RECT 19.37 57.79 19.53 67.9 ;
      RECT 18.81 6.24 19.41 6.84 ;
      RECT 19.01 56.99 19.41 57.29 ;
      RECT 19.21 48.24 19.37 50.5 ;
      RECT 19.14 26.68 19.3 28.17 ;
      RECT 19.13 29.97 19.29 34.08 ;
      RECT 19.13 39.34 19.29 43.45 ;
      RECT 18.89 57.79 19.05 62.72 ;
      RECT 18.65 29.97 18.81 32.28 ;
      RECT 18.65 35.23 18.81 36.31 ;
      RECT 18.65 37.11 18.81 38.19 ;
      RECT 18.65 41.14 18.81 43.45 ;
      RECT 18.45 12.28 18.77 12.76 ;
      RECT 18.25 8.96 18.76 9.17 ;
      RECT 18.57 21.73 18.73 22.33 ;
      RECT 18.57 22.49 18.73 23.06 ;
      RECT 18.41 57.79 18.57 62.72 ;
      RECT 18.27 15.09 18.55 15.41 ;
      RECT 17.01 6.24 18.41 6.84 ;
      RECT 18.25 47.88 18.41 51.16 ;
      RECT 17.91 36.21 18.11 36.95 ;
      RECT 17.93 21.45 18.09 24.52 ;
      RECT 17.93 29.32 18.09 34.08 ;
      RECT 17.93 39.34 18.09 46.59 ;
      RECT 17.93 47.59 18.09 51.92 ;
      RECT 17.93 52.64 18.09 56.5 ;
      RECT 17.61 47.83 17.77 51.16 ;
      RECT 17.45 57.79 17.61 62.72 ;
      RECT 17.21 29.97 17.37 32.28 ;
      RECT 17.21 35.23 17.37 36.31 ;
      RECT 17.21 37.11 17.37 38.19 ;
      RECT 17.21 41.14 17.37 43.45 ;
      RECT 9.29 15.46 17.13 16.9 ;
      RECT 16.97 57.79 17.13 62.72 ;
      RECT 16.61 56.99 17.01 57.29 ;
      RECT 16.73 29.97 16.89 34.08 ;
      RECT 16.73 39.34 16.89 43.45 ;
      RECT 16.65 48.24 16.81 50.5 ;
      RECT 16.49 57.79 16.65 67.9 ;
      RECT 14.61 510.54 16.61 510.94 ;
      RECT 14.61 6.24 16.59 6.84 ;
      RECT 16.25 29.97 16.41 32.28 ;
      RECT 16.25 35.23 16.41 36.31 ;
      RECT 16.25 37.11 16.41 38.19 ;
      RECT 16.25 41.14 16.41 43.45 ;
      RECT 10.19 21.67 16.23 21.95 ;
      RECT 15.51 36.21 15.71 36.95 ;
      RECT 15.53 29.32 15.69 34.08 ;
      RECT 15.53 39.34 15.69 46.59 ;
      RECT 15.53 47.59 15.69 51.11 ;
      RECT 15.53 51.34 15.69 53.67 ;
      RECT 15.53 54.16 15.69 56.5 ;
      RECT 14.81 29.97 14.97 32.28 ;
      RECT 14.81 35.23 14.97 36.31 ;
      RECT 14.81 37.11 14.97 38.19 ;
      RECT 14.81 41.14 14.97 43.45 ;
      RECT 14.57 57.79 14.73 67.9 ;
      RECT 14.21 56.99 14.61 57.29 ;
      RECT 14.41 48.24 14.57 50.5 ;
      RECT 14.33 29.97 14.49 34.08 ;
      RECT 14.33 39.34 14.49 43.45 ;
      RECT 14.09 57.79 14.25 62.72 ;
      RECT 12.21 6.24 14.19 6.84 ;
      RECT 13.85 29.97 14.01 32.28 ;
      RECT 13.85 35.23 14.01 36.31 ;
      RECT 13.85 37.11 14.01 38.19 ;
      RECT 13.85 41.14 14.01 43.45 ;
      RECT 13.61 57.79 13.77 62.72 ;
      RECT 13.45 47.88 13.61 51.16 ;
      RECT 12.93 9.36 13.49 9.52 ;
      RECT 12.93 11.3 13.49 11.46 ;
      RECT 12.93 14.68 13.49 14.84 ;
      RECT 12.93 19.63 13.49 19.79 ;
      RECT 13.11 36.21 13.31 36.95 ;
      RECT 13.13 29.32 13.29 34.08 ;
      RECT 13.13 39.34 13.29 46.59 ;
      RECT 13.13 47.59 13.29 51.92 ;
      RECT 13.13 52.64 13.29 56.5 ;
      RECT 12.81 47.88 12.97 51.16 ;
      RECT 12.65 57.79 12.81 62.72 ;
      RECT 12.41 29.97 12.57 32.28 ;
      RECT 12.41 35.23 12.57 36.31 ;
      RECT 12.41 37.11 12.57 38.19 ;
      RECT 12.41 41.14 12.57 43.45 ;
      RECT 12.17 57.79 12.33 62.72 ;
      RECT 11.81 56.99 12.21 57.29 ;
      RECT 11.93 29.97 12.09 34.08 ;
      RECT 11.93 39.34 12.09 43.45 ;
      RECT 11.85 48.24 12.01 50.5 ;
      RECT 11.69 57.79 11.85 67.9 ;
      RECT 9.81 510.54 11.81 510.94 ;
      RECT 9.81 6.24 11.79 6.84 ;
      RECT 11.45 29.97 11.61 32.28 ;
      RECT 11.45 35.23 11.61 36.31 ;
      RECT 11.45 37.11 11.61 38.19 ;
      RECT 11.45 41.14 11.61 43.45 ;
      RECT 10.71 36.21 10.91 36.95 ;
      RECT 10.73 29.32 10.89 34.08 ;
      RECT 10.73 39.34 10.89 46.59 ;
      RECT 10.73 47.59 10.89 51.11 ;
      RECT 10.73 51.34 10.89 53.67 ;
      RECT 10.73 54.16 10.89 56.5 ;
      RECT 10.01 29.97 10.17 32.28 ;
      RECT 10.01 35.23 10.17 36.31 ;
      RECT 10.01 37.11 10.17 38.19 ;
      RECT 10.01 41.14 10.17 43.45 ;
      RECT 9.77 57.79 9.93 67.9 ;
      RECT 9.41 56.99 9.81 57.29 ;
      RECT 9.61 48.24 9.77 50.5 ;
      RECT 9.53 29.97 9.69 34.08 ;
      RECT 9.53 39.34 9.69 43.45 ;
      RECT 9.29 57.79 9.45 62.72 ;
      RECT 7.41 6.24 9.41 6.84 ;
      RECT 9.05 29.97 9.21 32.28 ;
      RECT 9.05 35.23 9.21 36.31 ;
      RECT 9.05 37.11 9.21 38.19 ;
      RECT 9.05 41.14 9.21 43.45 ;
      RECT 8.81 57.79 8.97 62.72 ;
      RECT 8.65 47.88 8.81 51.16 ;
      RECT 8.31 36.21 8.51 36.95 ;
      RECT 8.33 29.32 8.49 34.08 ;
      RECT 8.33 39.34 8.49 46.59 ;
      RECT 8.33 47.59 8.49 51.92 ;
      RECT 8.33 52.64 8.49 56.5 ;
      RECT 6.75 10.92 7.03 11.4 ;
      RECT 6.75 18.87 7.03 19.35 ;
      RECT 6.75 14.87 7.02 15.29 ;
      RECT 6.75 9.34 7 9.78 ;
      RECT 6.24 7.94 6.82 9.14 ;
      RECT 6.24 17.26 6.82 18.46 ;
      RECT 6.24 25.81 6.82 27.81 ;
      RECT 6.24 35.91 6.82 36.91 ;
      RECT 6.24 50.24 6.82 51.24 ;
      RECT 6.24 57.02 6.82 58.02 ;
      RECT 6.24 60.6 6.82 61.6 ;
      RECT 6.24 62.45 6.82 63.45 ;
      RECT 6.24 69.16 6.82 69.96 ;
      RECT 6.24 72.56 6.82 73.36 ;
      RECT 6.24 75.96 6.82 76.76 ;
      RECT 6.24 79.36 6.82 80.16 ;
      RECT 6.24 82.76 6.82 83.56 ;
      RECT 6.24 86.16 6.82 86.96 ;
      RECT 6.24 89.56 6.82 90.36 ;
      RECT 6.24 92.96 6.82 93.76 ;
      RECT 6.24 96.36 6.82 97.16 ;
      RECT 6.24 99.76 6.82 100.56 ;
      RECT 6.24 103.16 6.82 103.96 ;
      RECT 6.24 106.56 6.82 107.36 ;
      RECT 6.24 109.96 6.82 110.76 ;
      RECT 6.24 113.36 6.82 114.16 ;
      RECT 6.24 116.76 6.82 117.56 ;
      RECT 6.24 120.16 6.82 120.96 ;
      RECT 6.24 123.56 6.82 124.36 ;
      RECT 6.24 126.96 6.82 127.76 ;
      RECT 6.24 130.36 6.82 131.16 ;
      RECT 6.24 133.76 6.82 134.56 ;
      RECT 6.24 137.16 6.82 137.96 ;
      RECT 6.24 140.56 6.82 141.36 ;
      RECT 6.24 143.96 6.82 144.76 ;
      RECT 6.24 147.36 6.82 148.16 ;
      RECT 6.24 150.76 6.82 151.56 ;
      RECT 6.24 154.16 6.82 154.96 ;
      RECT 6.24 157.56 6.82 158.36 ;
      RECT 6.24 160.96 6.82 161.76 ;
      RECT 6.24 164.36 6.82 165.16 ;
      RECT 6.24 167.76 6.82 168.56 ;
      RECT 6.24 171.16 6.82 171.96 ;
      RECT 6.24 174.56 6.82 175.36 ;
      RECT 6.24 177.96 6.82 178.76 ;
      RECT 6.24 181.36 6.82 182.16 ;
      RECT 6.24 184.76 6.82 185.56 ;
      RECT 6.24 188.16 6.82 188.96 ;
      RECT 6.24 191.56 6.82 192.36 ;
      RECT 6.24 194.96 6.82 195.76 ;
      RECT 6.24 198.36 6.82 199.16 ;
      RECT 6.24 201.76 6.82 202.56 ;
      RECT 6.24 205.16 6.82 205.96 ;
      RECT 6.24 208.56 6.82 209.36 ;
      RECT 6.24 211.96 6.82 212.76 ;
      RECT 6.24 215.36 6.82 216.16 ;
      RECT 6.24 218.76 6.82 219.56 ;
      RECT 6.24 222.16 6.82 222.96 ;
      RECT 6.24 225.56 6.82 226.36 ;
      RECT 6.24 228.96 6.82 229.76 ;
      RECT 6.24 232.36 6.82 233.16 ;
      RECT 6.24 235.76 6.82 236.56 ;
      RECT 6.24 239.16 6.82 239.96 ;
      RECT 6.24 242.56 6.82 243.36 ;
      RECT 6.24 245.96 6.82 246.76 ;
      RECT 6.24 249.36 6.82 250.16 ;
      RECT 6.24 252.76 6.82 253.56 ;
      RECT 6.24 256.16 6.82 256.96 ;
      RECT 6.24 259.56 6.82 260.36 ;
      RECT 6.24 262.96 6.82 263.76 ;
      RECT 6.24 266.36 6.82 267.16 ;
      RECT 6.24 269.76 6.82 270.56 ;
      RECT 6.24 273.16 6.82 273.96 ;
      RECT 6.24 276.56 6.82 277.36 ;
      RECT 6.24 279.96 6.82 280.76 ;
      RECT 6.24 283.36 6.82 284.16 ;
      RECT 6.24 286.76 6.82 287.56 ;
      RECT 6.24 290.16 6.82 290.96 ;
      RECT 6.24 293.56 6.82 294.36 ;
      RECT 6.24 296.96 6.82 297.76 ;
      RECT 6.24 300.36 6.82 301.16 ;
      RECT 6.24 303.76 6.82 304.56 ;
      RECT 6.24 307.16 6.82 307.96 ;
      RECT 6.24 310.56 6.82 311.36 ;
      RECT 6.24 313.96 6.82 314.76 ;
      RECT 6.24 317.36 6.82 318.16 ;
      RECT 6.24 320.76 6.82 321.56 ;
      RECT 6.24 324.16 6.82 324.96 ;
      RECT 6.24 327.56 6.82 328.36 ;
      RECT 6.24 330.96 6.82 331.76 ;
      RECT 6.24 334.36 6.82 335.16 ;
      RECT 6.24 337.76 6.82 338.56 ;
      RECT 6.24 341.16 6.82 341.96 ;
      RECT 6.24 344.56 6.82 345.36 ;
      RECT 6.24 347.96 6.82 348.76 ;
      RECT 6.24 351.36 6.82 352.16 ;
      RECT 6.24 354.76 6.82 355.56 ;
      RECT 6.24 358.16 6.82 358.96 ;
      RECT 6.24 361.56 6.82 362.36 ;
      RECT 6.24 364.96 6.82 365.76 ;
      RECT 6.24 368.36 6.82 369.16 ;
      RECT 6.24 371.76 6.82 372.56 ;
      RECT 6.24 375.16 6.82 375.96 ;
      RECT 6.24 378.56 6.82 379.36 ;
      RECT 6.24 381.96 6.82 382.76 ;
      RECT 6.24 385.36 6.82 386.16 ;
      RECT 6.24 388.76 6.82 389.56 ;
      RECT 6.24 392.16 6.82 392.96 ;
      RECT 6.24 395.56 6.82 396.36 ;
      RECT 6.24 398.96 6.82 399.76 ;
      RECT 6.24 402.36 6.82 403.16 ;
      RECT 6.24 405.76 6.82 406.56 ;
      RECT 6.24 409.16 6.82 409.96 ;
      RECT 6.24 412.56 6.82 413.36 ;
      RECT 6.24 415.96 6.82 416.76 ;
      RECT 6.24 419.36 6.82 420.16 ;
      RECT 6.24 422.76 6.82 423.56 ;
      RECT 6.24 426.16 6.82 426.96 ;
      RECT 6.24 429.56 6.82 430.36 ;
      RECT 6.24 432.96 6.82 433.76 ;
      RECT 6.24 436.36 6.82 437.16 ;
      RECT 6.24 439.76 6.82 440.56 ;
      RECT 6.24 443.16 6.82 443.96 ;
      RECT 6.24 446.56 6.82 447.36 ;
      RECT 6.24 449.96 6.82 450.76 ;
      RECT 6.24 453.36 6.82 454.16 ;
      RECT 6.24 456.76 6.82 457.56 ;
      RECT 6.24 460.16 6.82 460.96 ;
      RECT 6.24 463.56 6.82 464.36 ;
      RECT 6.24 466.96 6.82 467.76 ;
      RECT 6.24 470.36 6.82 471.16 ;
      RECT 6.24 473.76 6.82 474.56 ;
      RECT 6.24 477.16 6.82 477.96 ;
      RECT 6.24 480.56 6.82 481.36 ;
      RECT 6.24 483.96 6.82 484.76 ;
      RECT 6.24 487.36 6.82 488.16 ;
      RECT 6.24 490.76 6.82 491.56 ;
      RECT 6.24 494.16 6.82 494.96 ;
      RECT 6.24 497.56 6.82 498.36 ;
      RECT 6.24 500.96 6.82 501.76 ;
      RECT 6.24 504.36 6.82 505.16 ;
      RECT 6.24 505.6 6.82 506 ;
      RECT 6.24 509 6.82 509.8 ;
    LAYER M2 ;
      RECT 233.76 7.94 234.36 9.14 ;
      RECT 222.49 8.34 222.69 9.14 ;
      RECT 203.29 8.34 203.49 9.14 ;
      RECT 182.89 8.34 183.09 9.14 ;
      RECT 163.69 8.34 163.89 9.14 ;
      RECT 76.71 8.34 76.91 9.14 ;
      RECT 57.51 8.34 57.71 9.14 ;
      RECT 37.11 8.34 37.31 9.14 ;
      RECT 17.91 8.34 18.11 9.14 ;
      RECT 6.24 7.94 6.84 9.14 ;
      RECT 6.24 8.34 234.36 8.74 ;
      RECT 88.61 17.66 151.71 19.86 ;
      RECT 233.76 17.26 234.36 18.46 ;
      RECT 6.24 17.26 6.84 18.46 ;
      RECT 6.24 17.66 234.36 18.06 ;
      RECT 233.36 21.41 234.36 22.21 ;
      RECT 6.24 21.41 7.24 22.21 ;
      RECT 6.24 21.71 234.36 22.11 ;
      RECT 222.49 21.41 234.36 22.11 ;
      RECT 212.89 21.41 213.09 22.11 ;
      RECT 182.89 21.41 203.49 22.11 ;
      RECT 173.29 21.41 173.49 22.11 ;
      RECT 76.71 21.41 163.89 22.11 ;
      RECT 67.11 21.41 67.31 22.11 ;
      RECT 37.11 21.41 57.71 22.11 ;
      RECT 27.51 21.41 27.71 22.11 ;
      RECT 6.24 21.41 18.11 22.11 ;
      RECT 233.36 25.81 234.36 27.81 ;
      RECT 6.24 25.81 7.24 27.81 ;
      RECT 6.24 26.91 234.36 27.31 ;
      RECT 219.41 26.31 234.36 27.31 ;
      RECT 209.81 26.11 216.17 27.31 ;
      RECT 215.97 25.48 216.17 27.31 ;
      RECT 179.81 26.31 206.57 27.31 ;
      RECT 206.37 25.48 206.57 27.31 ;
      RECT 170.21 26.11 176.57 27.31 ;
      RECT 176.37 25.48 176.57 27.31 ;
      RECT 73.63 26.31 166.97 27.31 ;
      RECT 166.77 25.48 166.97 27.31 ;
      RECT 64.03 26.11 70.39 27.31 ;
      RECT 70.19 25.48 70.39 27.31 ;
      RECT 34.03 26.31 60.79 27.31 ;
      RECT 60.59 25.48 60.79 27.31 ;
      RECT 24.43 26.11 30.79 27.31 ;
      RECT 30.59 25.48 30.79 27.31 ;
      RECT 6.24 26.31 21.19 27.31 ;
      RECT 20.99 25.48 21.19 27.31 ;
      RECT 219.41 26.11 222.59 27.31 ;
      RECT 203.39 26.11 206.57 27.31 ;
      RECT 179.81 26.11 182.99 27.31 ;
      RECT 163.79 26.11 166.97 27.31 ;
      RECT 73.63 26.11 76.81 27.31 ;
      RECT 57.61 26.11 60.79 27.31 ;
      RECT 34.03 26.11 37.21 27.31 ;
      RECT 18.01 26.11 21.19 27.31 ;
      RECT 219.41 25.48 219.61 27.31 ;
      RECT 209.81 25.48 210.01 27.31 ;
      RECT 179.81 25.48 180.01 27.31 ;
      RECT 170.21 25.48 170.41 27.31 ;
      RECT 73.63 25.48 73.83 27.31 ;
      RECT 64.03 25.48 64.23 27.31 ;
      RECT 34.03 25.48 34.23 27.31 ;
      RECT 24.43 25.48 24.63 27.31 ;
      RECT 85.81 35.75 87.01 35.95 ;
      RECT 86.81 32.98 87.01 35.95 ;
      RECT 85.81 34.65 87.01 34.85 ;
      RECT 6.24 32.98 234.36 33.98 ;
      RECT 6.24 36.25 234.36 36.91 ;
      RECT 233.76 35.91 234.36 36.91 ;
      RECT 87.81 35.91 153.54 36.91 ;
      RECT 6.24 35.91 6.84 36.91 ;
      RECT 6.24 39.44 234.36 40.44 ;
      RECT 138.92 37.58 139.12 40.44 ;
      RECT 137 37.58 137.2 40.44 ;
      RECT 89.4 39.17 95.02 40.44 ;
      RECT 94.82 37.58 95.02 40.44 ;
      RECT 86.81 37.21 87.01 40.44 ;
      RECT 89.4 37.58 89.6 40.44 ;
      RECT 85.81 38.81 87.01 39.01 ;
      RECT 85.81 37.21 87.01 37.41 ;
      RECT 152.09 62.45 234.36 63.45 ;
      RECT 6.24 62.45 87.61 63.45 ;
      RECT 86.61 60.6 87.61 63.45 ;
      RECT 152.09 60.6 153.09 63.45 ;
      RECT 6.24 60.6 234.36 61.6 ;
      RECT 232.39 510.34 233.19 510.94 ;
      RECT 231.19 510.34 231.99 510.94 ;
      RECT 231.19 510.34 233.39 510.74 ;
      RECT 233.09 68.04 233.29 510.74 ;
      RECT 232.29 68.04 232.49 510.74 ;
      RECT 231.49 65.96 231.69 510.94 ;
      RECT 233.09 506.6 234.36 508.6 ;
      RECT 233.09 502.66 234.36 503.46 ;
      RECT 233.09 499.26 234.36 500.06 ;
      RECT 233.09 495.86 234.36 496.66 ;
      RECT 233.09 492.46 234.36 493.26 ;
      RECT 233.09 489.06 234.36 489.86 ;
      RECT 233.09 485.66 234.36 486.46 ;
      RECT 233.09 482.26 234.36 483.06 ;
      RECT 233.09 478.86 234.36 479.66 ;
      RECT 233.09 475.46 234.36 476.26 ;
      RECT 233.09 472.06 234.36 472.86 ;
      RECT 233.09 468.66 234.36 469.46 ;
      RECT 233.09 465.26 234.36 466.06 ;
      RECT 233.09 461.86 234.36 462.66 ;
      RECT 233.09 458.46 234.36 459.26 ;
      RECT 233.09 455.06 234.36 455.86 ;
      RECT 233.09 451.66 234.36 452.46 ;
      RECT 233.09 448.26 234.36 449.06 ;
      RECT 233.09 444.86 234.36 445.66 ;
      RECT 233.09 441.46 234.36 442.26 ;
      RECT 233.09 438.06 234.36 438.86 ;
      RECT 233.09 434.66 234.36 435.46 ;
      RECT 233.09 431.26 234.36 432.06 ;
      RECT 233.09 427.86 234.36 428.66 ;
      RECT 233.09 424.46 234.36 425.26 ;
      RECT 233.09 421.06 234.36 421.86 ;
      RECT 233.09 417.66 234.36 418.46 ;
      RECT 233.09 414.26 234.36 415.06 ;
      RECT 233.09 410.86 234.36 411.66 ;
      RECT 233.09 407.46 234.36 408.26 ;
      RECT 233.09 404.06 234.36 404.86 ;
      RECT 233.09 400.66 234.36 401.46 ;
      RECT 233.09 397.26 234.36 398.06 ;
      RECT 233.09 393.86 234.36 394.66 ;
      RECT 233.09 390.46 234.36 391.26 ;
      RECT 233.09 387.06 234.36 387.86 ;
      RECT 233.09 383.66 234.36 384.46 ;
      RECT 233.09 380.26 234.36 381.06 ;
      RECT 233.09 376.86 234.36 377.66 ;
      RECT 233.09 373.46 234.36 374.26 ;
      RECT 233.09 370.06 234.36 370.86 ;
      RECT 233.09 366.66 234.36 367.46 ;
      RECT 233.09 363.26 234.36 364.06 ;
      RECT 233.09 359.86 234.36 360.66 ;
      RECT 233.09 356.46 234.36 357.26 ;
      RECT 233.09 353.06 234.36 353.86 ;
      RECT 233.09 349.66 234.36 350.46 ;
      RECT 233.09 346.26 234.36 347.06 ;
      RECT 233.09 342.86 234.36 343.66 ;
      RECT 233.09 339.46 234.36 340.26 ;
      RECT 233.09 336.06 234.36 336.86 ;
      RECT 233.09 332.66 234.36 333.46 ;
      RECT 233.09 329.26 234.36 330.06 ;
      RECT 233.09 325.86 234.36 326.66 ;
      RECT 233.09 322.46 234.36 323.26 ;
      RECT 233.09 319.06 234.36 319.86 ;
      RECT 233.09 315.66 234.36 316.46 ;
      RECT 233.09 312.26 234.36 313.06 ;
      RECT 233.09 308.86 234.36 309.66 ;
      RECT 233.09 305.46 234.36 306.26 ;
      RECT 233.09 302.06 234.36 302.86 ;
      RECT 233.09 298.66 234.36 299.46 ;
      RECT 233.09 295.26 234.36 296.06 ;
      RECT 233.09 291.86 234.36 292.66 ;
      RECT 233.09 288.46 234.36 289.26 ;
      RECT 233.09 285.06 234.36 285.86 ;
      RECT 233.09 281.66 234.36 282.46 ;
      RECT 233.09 278.26 234.36 279.06 ;
      RECT 233.09 274.86 234.36 275.66 ;
      RECT 233.09 271.46 234.36 272.26 ;
      RECT 233.09 268.06 234.36 268.86 ;
      RECT 233.09 264.66 234.36 265.46 ;
      RECT 233.09 261.26 234.36 262.06 ;
      RECT 233.09 257.86 234.36 258.66 ;
      RECT 233.09 254.46 234.36 255.26 ;
      RECT 233.09 251.06 234.36 251.86 ;
      RECT 233.09 247.66 234.36 248.46 ;
      RECT 233.09 244.26 234.36 245.06 ;
      RECT 233.09 240.86 234.36 241.66 ;
      RECT 233.09 237.46 234.36 238.26 ;
      RECT 233.09 234.06 234.36 234.86 ;
      RECT 233.09 230.66 234.36 231.46 ;
      RECT 233.09 227.26 234.36 228.06 ;
      RECT 233.09 223.86 234.36 224.66 ;
      RECT 233.09 220.46 234.36 221.26 ;
      RECT 233.09 217.06 234.36 217.86 ;
      RECT 233.09 213.66 234.36 214.46 ;
      RECT 233.09 210.26 234.36 211.06 ;
      RECT 233.09 206.86 234.36 207.66 ;
      RECT 233.09 203.46 234.36 204.26 ;
      RECT 233.09 200.06 234.36 200.86 ;
      RECT 233.09 196.66 234.36 197.46 ;
      RECT 233.09 193.26 234.36 194.06 ;
      RECT 233.09 189.86 234.36 190.66 ;
      RECT 233.09 186.46 234.36 187.26 ;
      RECT 233.09 183.06 234.36 183.86 ;
      RECT 233.09 179.66 234.36 180.46 ;
      RECT 233.09 176.26 234.36 177.06 ;
      RECT 233.09 172.86 234.36 173.66 ;
      RECT 233.09 169.46 234.36 170.26 ;
      RECT 233.09 166.06 234.36 166.86 ;
      RECT 233.09 162.66 234.36 163.46 ;
      RECT 233.09 159.26 234.36 160.06 ;
      RECT 233.09 155.86 234.36 156.66 ;
      RECT 233.09 152.46 234.36 153.26 ;
      RECT 233.09 149.06 234.36 149.86 ;
      RECT 233.09 145.66 234.36 146.46 ;
      RECT 233.09 142.26 234.36 143.06 ;
      RECT 233.09 138.86 234.36 139.66 ;
      RECT 233.09 135.46 234.36 136.26 ;
      RECT 233.09 132.06 234.36 132.86 ;
      RECT 233.09 128.66 234.36 129.46 ;
      RECT 233.09 125.26 234.36 126.06 ;
      RECT 233.09 121.86 234.36 122.66 ;
      RECT 233.09 118.46 234.36 119.26 ;
      RECT 233.09 115.06 234.36 115.86 ;
      RECT 233.09 111.66 234.36 112.46 ;
      RECT 233.09 108.26 234.36 109.06 ;
      RECT 233.09 104.86 234.36 105.66 ;
      RECT 233.09 101.46 234.36 102.26 ;
      RECT 233.09 98.06 234.36 98.86 ;
      RECT 233.09 94.66 234.36 95.46 ;
      RECT 233.09 91.26 234.36 92.06 ;
      RECT 233.09 87.86 234.36 88.66 ;
      RECT 233.09 84.46 234.36 85.26 ;
      RECT 233.09 81.06 234.36 81.86 ;
      RECT 233.09 77.66 234.36 78.46 ;
      RECT 233.09 74.26 234.36 75.06 ;
      RECT 233.09 70.86 234.36 71.66 ;
      RECT 232.29 68.04 233.29 68.24 ;
      RECT 152.09 10.98 232.39 11.78 ;
      RECT 152.09 10.98 233.76 11.34 ;
      RECT 222.09 14.34 222.29 15.4 ;
      RECT 203.69 14.34 203.89 15.4 ;
      RECT 182.49 14.34 182.69 15.4 ;
      RECT 164.09 14.34 164.29 15.4 ;
      RECT 76.31 14.34 76.51 15.4 ;
      RECT 57.91 14.34 58.11 15.4 ;
      RECT 36.71 14.34 36.91 15.4 ;
      RECT 18.31 14.34 18.51 15.4 ;
      RECT 6.84 14.98 233.76 15.18 ;
      RECT 150.62 14.34 233.76 15.18 ;
      RECT 142.15 14.35 233.76 15.18 ;
      RECT 6.84 14.34 87.18 15.18 ;
      RECT 87.63 14.35 233.76 14.78 ;
      RECT 231.59 35.75 233.36 35.95 ;
      RECT 233.14 34.65 233.36 35.95 ;
      RECT 231.59 34.65 233.36 34.85 ;
      RECT 231.59 38.81 233.36 39.01 ;
      RECT 233.14 37.21 233.36 39.01 ;
      RECT 231.59 37.21 233.36 37.41 ;
      RECT 231.89 65.25 232.09 505.18 ;
      RECT 231.49 65.25 232.09 65.45 ;
      RECT 231.49 63.99 231.69 65.45 ;
      RECT 231.61 58.57 231.81 59.17 ;
      RECT 230.29 58.57 230.49 59.17 ;
      RECT 230.29 58.57 231.81 58.77 ;
      RECT 231.49 37.91 231.69 38.61 ;
      RECT 231.29 37.91 231.69 38.11 ;
      RECT 212.39 38.81 231.09 39.01 ;
      RECT 230.89 37.61 231.09 39.01 ;
      RECT 228.49 37.61 228.69 39.01 ;
      RECT 226.09 37.61 226.29 39.01 ;
      RECT 223.69 37.61 223.89 39.01 ;
      RECT 221.29 37.61 221.49 39.01 ;
      RECT 218.89 37.61 219.09 39.01 ;
      RECT 216.49 37.61 216.69 39.01 ;
      RECT 214.09 37.61 214.29 39.01 ;
      RECT 229.89 63.99 230.09 505.18 ;
      RECT 230.69 63.99 230.89 65.05 ;
      RECT 229.89 63.99 230.89 64.19 ;
      RECT 230.69 65.25 230.89 505.18 ;
      RECT 230.29 65.25 230.89 65.45 ;
      RECT 230.29 64.39 230.49 65.45 ;
      RECT 228.79 510.34 230.79 510.94 ;
      RECT 230.29 65.96 230.49 510.94 ;
      RECT 230.29 37.91 230.49 38.61 ;
      RECT 230.29 37.91 230.69 38.11 ;
      RECT 229.49 63.99 229.69 505.18 ;
      RECT 228.69 63.99 228.89 65.05 ;
      RECT 228.69 63.99 229.69 64.19 ;
      RECT 229.09 37.91 229.29 38.61 ;
      RECT 228.89 37.91 229.29 38.11 ;
      RECT 229.09 58.57 229.29 59.17 ;
      RECT 227.77 58.57 227.97 59.17 ;
      RECT 227.77 58.57 229.29 58.77 ;
      RECT 228.69 65.25 228.89 505.18 ;
      RECT 228.69 65.25 229.29 65.45 ;
      RECT 229.09 64.39 229.29 65.45 ;
      RECT 227.59 510.34 228.39 510.94 ;
      RECT 226.39 510.34 227.19 510.94 ;
      RECT 226.39 510.34 228.39 510.74 ;
      RECT 226.69 65.96 226.89 510.94 ;
      RECT 227.89 37.91 228.09 38.61 ;
      RECT 227.89 37.91 228.29 38.11 ;
      RECT 227.49 65.25 227.69 505.18 ;
      RECT 227.49 65.25 228.09 65.45 ;
      RECT 227.89 63.99 228.09 65.45 ;
      RECT 227.09 65.25 227.29 505.18 ;
      RECT 226.69 65.25 227.29 65.45 ;
      RECT 226.69 63.99 226.89 65.45 ;
      RECT 226.81 58.57 227.01 59.17 ;
      RECT 225.49 58.57 225.69 59.17 ;
      RECT 225.49 58.57 227.01 58.77 ;
      RECT 226.69 37.91 226.89 38.61 ;
      RECT 226.49 37.91 226.89 38.11 ;
      RECT 225.09 63.99 225.29 505.18 ;
      RECT 225.89 63.99 226.09 65.05 ;
      RECT 225.09 63.99 226.09 64.19 ;
      RECT 225.89 65.25 226.09 505.18 ;
      RECT 225.49 65.25 226.09 65.45 ;
      RECT 225.49 64.39 225.69 65.45 ;
      RECT 223.99 510.34 225.99 510.94 ;
      RECT 225.49 65.96 225.69 510.94 ;
      RECT 225.49 37.91 225.69 38.61 ;
      RECT 225.49 37.91 225.89 38.11 ;
      RECT 224.69 63.99 224.89 505.18 ;
      RECT 223.89 63.99 224.09 65.05 ;
      RECT 223.89 63.99 224.89 64.19 ;
      RECT 224.29 37.91 224.49 38.61 ;
      RECT 224.09 37.91 224.49 38.11 ;
      RECT 224.29 58.57 224.49 59.17 ;
      RECT 222.97 58.57 223.17 59.17 ;
      RECT 222.97 58.57 224.49 58.77 ;
      RECT 223.89 65.25 224.09 505.18 ;
      RECT 223.89 65.25 224.49 65.45 ;
      RECT 224.29 64.39 224.49 65.45 ;
      RECT 222.79 510.34 223.59 510.94 ;
      RECT 221.59 510.34 222.39 510.94 ;
      RECT 221.59 510.34 223.59 510.74 ;
      RECT 221.89 65.96 222.09 510.94 ;
      RECT 223.09 37.91 223.29 38.61 ;
      RECT 223.09 37.91 223.49 38.11 ;
      RECT 222.69 65.25 222.89 505.18 ;
      RECT 222.69 65.25 223.29 65.45 ;
      RECT 223.09 63.99 223.29 65.45 ;
      RECT 222.29 65.25 222.49 505.18 ;
      RECT 221.89 65.25 222.49 65.45 ;
      RECT 221.89 63.99 222.09 65.45 ;
      RECT 222.01 58.57 222.21 59.17 ;
      RECT 220.69 58.57 220.89 59.17 ;
      RECT 220.69 58.57 222.21 58.77 ;
      RECT 220.13 24.85 222.19 25.05 ;
      RECT 221.99 24.22 222.19 25.05 ;
      RECT 215.31 12.98 218.99 13.18 ;
      RECT 218.79 12.58 218.99 13.18 ;
      RECT 218.79 12.58 222.09 12.78 ;
      RECT 221.89 37.91 222.09 38.61 ;
      RECT 221.69 37.91 222.09 38.11 ;
      RECT 219.67 23.59 222.05 23.79 ;
      RECT 221.85 22.77 222.05 23.79 ;
      RECT 217.69 22.71 217.89 26.71 ;
      RECT 214.11 22.71 221.47 22.91 ;
      RECT 220.29 63.99 220.49 505.18 ;
      RECT 221.09 63.99 221.29 65.05 ;
      RECT 220.29 63.99 221.29 64.19 ;
      RECT 221.09 65.25 221.29 505.18 ;
      RECT 220.69 65.25 221.29 65.45 ;
      RECT 220.69 64.39 220.89 65.45 ;
      RECT 219.19 510.34 221.19 510.94 ;
      RECT 220.69 65.96 220.89 510.94 ;
      RECT 220.69 37.91 220.89 38.61 ;
      RECT 220.69 37.91 221.09 38.11 ;
      RECT 219.89 63.99 220.09 505.18 ;
      RECT 219.09 63.99 219.29 65.05 ;
      RECT 219.09 63.99 220.09 64.19 ;
      RECT 214.49 16.9 220.06 17.1 ;
      RECT 219.38 15.79 219.58 17.1 ;
      RECT 218.83 15.79 219.58 15.99 ;
      RECT 219.49 37.91 219.69 38.61 ;
      RECT 219.29 37.91 219.69 38.11 ;
      RECT 219.49 58.57 219.69 59.17 ;
      RECT 218.17 58.57 218.37 59.17 ;
      RECT 218.17 58.57 219.69 58.77 ;
      RECT 219.09 65.25 219.29 505.18 ;
      RECT 219.09 65.25 219.69 65.45 ;
      RECT 219.49 64.39 219.69 65.45 ;
      RECT 217.45 16.27 219.18 16.47 ;
      RECT 214.03 16.1 217.65 16.3 ;
      RECT 218.09 23.11 218.29 26.31 ;
      RECT 218.09 23.11 218.89 23.31 ;
      RECT 218.49 26.46 218.89 26.66 ;
      RECT 218.49 24.68 218.69 26.66 ;
      RECT 217.99 510.34 218.79 510.94 ;
      RECT 216.79 510.34 217.59 510.94 ;
      RECT 216.79 510.34 218.79 510.74 ;
      RECT 217.09 65.96 217.29 510.94 ;
      RECT 218.29 37.91 218.49 38.61 ;
      RECT 218.29 37.91 218.69 38.11 ;
      RECT 217.89 65.25 218.09 505.18 ;
      RECT 217.89 65.25 218.49 65.45 ;
      RECT 218.29 63.99 218.49 65.45 ;
      RECT 217.49 65.25 217.69 505.18 ;
      RECT 217.09 65.25 217.69 65.45 ;
      RECT 217.09 63.99 217.29 65.45 ;
      RECT 217.29 23.11 217.49 26.31 ;
      RECT 216.69 23.11 217.49 23.31 ;
      RECT 217.21 58.57 217.41 59.17 ;
      RECT 215.89 58.57 216.09 59.17 ;
      RECT 215.89 58.57 217.41 58.77 ;
      RECT 217.09 37.91 217.29 38.61 ;
      RECT 216.89 37.91 217.29 38.11 ;
      RECT 216.69 26.46 217.09 26.66 ;
      RECT 216.89 24.68 217.09 26.66 ;
      RECT 215.49 63.99 215.69 505.18 ;
      RECT 216.29 63.99 216.49 65.05 ;
      RECT 215.49 63.99 216.49 64.19 ;
      RECT 216.29 65.25 216.49 505.18 ;
      RECT 215.89 65.25 216.49 65.45 ;
      RECT 215.89 64.39 216.09 65.45 ;
      RECT 214.39 510.34 216.39 510.94 ;
      RECT 215.89 65.96 216.09 510.94 ;
      RECT 215.89 37.91 216.09 38.61 ;
      RECT 215.89 37.91 216.29 38.11 ;
      RECT 213.53 23.59 215.91 23.79 ;
      RECT 213.53 22.77 213.73 23.79 ;
      RECT 213.39 24.85 215.45 25.05 ;
      RECT 213.39 24.22 213.59 25.05 ;
      RECT 215.09 63.99 215.29 505.18 ;
      RECT 214.29 63.99 214.49 65.05 ;
      RECT 214.29 63.99 215.29 64.19 ;
      RECT 214.99 15.38 215.19 15.9 ;
      RECT 214.49 15.38 215.19 15.58 ;
      RECT 214.69 37.91 214.89 38.61 ;
      RECT 214.49 37.91 214.89 38.11 ;
      RECT 214.69 58.57 214.89 59.17 ;
      RECT 213.37 58.57 213.57 59.17 ;
      RECT 213.37 58.57 214.89 58.77 ;
      RECT 214.29 65.25 214.49 505.18 ;
      RECT 214.29 65.25 214.89 65.45 ;
      RECT 214.69 64.39 214.89 65.45 ;
      RECT 213.19 510.34 213.99 510.94 ;
      RECT 211.99 510.34 212.79 510.94 ;
      RECT 211.99 510.34 213.99 510.74 ;
      RECT 212.29 65.96 212.49 510.94 ;
      RECT 213.49 37.91 213.69 38.61 ;
      RECT 213.49 37.91 213.89 38.11 ;
      RECT 213.09 65.25 213.29 505.18 ;
      RECT 213.09 65.25 213.69 65.45 ;
      RECT 213.49 63.99 213.69 65.45 ;
      RECT 212.69 65.25 212.89 505.18 ;
      RECT 212.29 65.25 212.89 65.45 ;
      RECT 212.29 63.99 212.49 65.45 ;
      RECT 212.41 58.57 212.61 59.17 ;
      RECT 211.09 58.57 211.29 59.17 ;
      RECT 211.09 58.57 212.61 58.77 ;
      RECT 210.53 24.85 212.59 25.05 ;
      RECT 212.39 24.22 212.59 25.05 ;
      RECT 212.29 37.91 212.49 38.61 ;
      RECT 212.09 37.91 212.49 38.11 ;
      RECT 210.07 23.59 212.45 23.79 ;
      RECT 212.25 22.77 212.45 23.79 ;
      RECT 206.8 16.27 208.53 16.47 ;
      RECT 208.33 16.1 211.95 16.3 ;
      RECT 191.99 38.81 211.89 39.01 ;
      RECT 211.69 37.61 211.89 39.01 ;
      RECT 209.29 37.61 209.49 39.01 ;
      RECT 206.89 37.61 207.09 39.01 ;
      RECT 204.49 37.61 204.69 39.01 ;
      RECT 202.09 37.61 202.29 39.01 ;
      RECT 199.69 37.61 199.89 39.01 ;
      RECT 197.29 37.61 197.49 39.01 ;
      RECT 194.89 37.61 195.09 39.01 ;
      RECT 208.09 22.71 208.29 26.71 ;
      RECT 204.51 22.71 211.87 22.91 ;
      RECT 210.69 63.99 210.89 505.18 ;
      RECT 211.49 63.99 211.69 65.05 ;
      RECT 210.69 63.99 211.69 64.19 ;
      RECT 211.49 65.25 211.69 505.18 ;
      RECT 211.09 65.25 211.69 65.45 ;
      RECT 211.09 64.39 211.29 65.45 ;
      RECT 209.59 510.34 211.59 510.94 ;
      RECT 211.09 65.96 211.29 510.94 ;
      RECT 210.79 15.38 210.99 15.9 ;
      RECT 210.79 15.38 211.49 15.58 ;
      RECT 205.92 16.9 211.49 17.1 ;
      RECT 206.4 15.79 206.6 17.1 ;
      RECT 206.4 15.79 207.15 15.99 ;
      RECT 211.09 37.91 211.29 38.61 ;
      RECT 211.09 37.91 211.49 38.11 ;
      RECT 206.99 12.98 210.67 13.18 ;
      RECT 206.99 12.58 207.19 13.18 ;
      RECT 203.89 12.58 207.19 12.78 ;
      RECT 210.29 63.99 210.49 505.18 ;
      RECT 209.49 63.99 209.69 65.05 ;
      RECT 209.49 63.99 210.49 64.19 ;
      RECT 209.89 37.91 210.09 38.61 ;
      RECT 209.69 37.91 210.09 38.11 ;
      RECT 209.89 58.57 210.09 59.17 ;
      RECT 208.57 58.57 208.77 59.17 ;
      RECT 208.57 58.57 210.09 58.77 ;
      RECT 209.49 65.25 209.69 505.18 ;
      RECT 209.49 65.25 210.09 65.45 ;
      RECT 209.89 64.39 210.09 65.45 ;
      RECT 208.49 23.11 208.69 26.31 ;
      RECT 208.49 23.11 209.29 23.31 ;
      RECT 208.89 26.46 209.29 26.66 ;
      RECT 208.89 24.68 209.09 26.66 ;
      RECT 208.39 510.34 209.19 510.94 ;
      RECT 207.19 510.34 207.99 510.94 ;
      RECT 207.19 510.34 209.19 510.74 ;
      RECT 207.49 65.96 207.69 510.94 ;
      RECT 208.69 37.91 208.89 38.61 ;
      RECT 208.69 37.91 209.09 38.11 ;
      RECT 208.29 65.25 208.49 505.18 ;
      RECT 208.29 65.25 208.89 65.45 ;
      RECT 208.69 63.99 208.89 65.45 ;
      RECT 207.89 65.25 208.09 505.18 ;
      RECT 207.49 65.25 208.09 65.45 ;
      RECT 207.49 63.99 207.69 65.45 ;
      RECT 207.69 23.11 207.89 26.31 ;
      RECT 207.09 23.11 207.89 23.31 ;
      RECT 207.61 58.57 207.81 59.17 ;
      RECT 206.29 58.57 206.49 59.17 ;
      RECT 206.29 58.57 207.81 58.77 ;
      RECT 207.49 37.91 207.69 38.61 ;
      RECT 207.29 37.91 207.69 38.11 ;
      RECT 207.09 26.46 207.49 26.66 ;
      RECT 207.29 24.68 207.49 26.66 ;
      RECT 205.89 63.99 206.09 505.18 ;
      RECT 206.69 63.99 206.89 65.05 ;
      RECT 205.89 63.99 206.89 64.19 ;
      RECT 206.69 65.25 206.89 505.18 ;
      RECT 206.29 65.25 206.89 65.45 ;
      RECT 206.29 64.39 206.49 65.45 ;
      RECT 204.79 510.34 206.79 510.94 ;
      RECT 206.29 65.96 206.49 510.94 ;
      RECT 206.29 37.91 206.49 38.61 ;
      RECT 206.29 37.91 206.69 38.11 ;
      RECT 203.93 23.59 206.31 23.79 ;
      RECT 203.93 22.77 204.13 23.79 ;
      RECT 203.79 24.85 205.85 25.05 ;
      RECT 203.79 24.22 203.99 25.05 ;
      RECT 205.49 63.99 205.69 505.18 ;
      RECT 204.69 63.99 204.89 65.05 ;
      RECT 204.69 63.99 205.69 64.19 ;
      RECT 205.09 37.91 205.29 38.61 ;
      RECT 204.89 37.91 205.29 38.11 ;
      RECT 205.09 58.57 205.29 59.17 ;
      RECT 203.77 58.57 203.97 59.17 ;
      RECT 203.77 58.57 205.29 58.77 ;
      RECT 204.69 65.25 204.89 505.18 ;
      RECT 204.69 65.25 205.29 65.45 ;
      RECT 205.09 64.39 205.29 65.45 ;
      RECT 203.59 510.34 204.39 510.94 ;
      RECT 202.39 510.34 203.19 510.94 ;
      RECT 202.39 510.34 204.39 510.74 ;
      RECT 202.69 65.96 202.89 510.94 ;
      RECT 203.89 37.91 204.09 38.61 ;
      RECT 203.89 37.91 204.29 38.11 ;
      RECT 203.49 65.25 203.69 505.18 ;
      RECT 203.49 65.25 204.09 65.45 ;
      RECT 203.89 63.99 204.09 65.45 ;
      RECT 203.09 65.25 203.29 505.18 ;
      RECT 202.69 65.25 203.29 65.45 ;
      RECT 202.69 63.99 202.89 65.45 ;
      RECT 202.81 58.57 203.01 59.17 ;
      RECT 201.49 58.57 201.69 59.17 ;
      RECT 201.49 58.57 203.01 58.77 ;
      RECT 202.69 37.91 202.89 38.61 ;
      RECT 202.49 37.91 202.89 38.11 ;
      RECT 201.09 63.99 201.29 505.18 ;
      RECT 201.89 63.99 202.09 65.05 ;
      RECT 201.09 63.99 202.09 64.19 ;
      RECT 201.89 65.25 202.09 505.18 ;
      RECT 201.49 65.25 202.09 65.45 ;
      RECT 201.49 64.39 201.69 65.45 ;
      RECT 199.99 510.34 201.99 510.94 ;
      RECT 201.49 65.96 201.69 510.94 ;
      RECT 201.49 37.91 201.69 38.61 ;
      RECT 201.49 37.91 201.89 38.11 ;
      RECT 200.69 63.99 200.89 505.18 ;
      RECT 199.89 63.99 200.09 65.05 ;
      RECT 199.89 63.99 200.89 64.19 ;
      RECT 200.29 37.91 200.49 38.61 ;
      RECT 200.09 37.91 200.49 38.11 ;
      RECT 200.29 58.57 200.49 59.17 ;
      RECT 198.97 58.57 199.17 59.17 ;
      RECT 198.97 58.57 200.49 58.77 ;
      RECT 199.89 65.25 200.09 505.18 ;
      RECT 199.89 65.25 200.49 65.45 ;
      RECT 200.29 64.39 200.49 65.45 ;
      RECT 198.79 510.34 199.59 510.94 ;
      RECT 197.59 510.34 198.39 510.94 ;
      RECT 197.59 510.34 199.59 510.74 ;
      RECT 197.89 65.96 198.09 510.94 ;
      RECT 199.09 37.91 199.29 38.61 ;
      RECT 199.09 37.91 199.49 38.11 ;
      RECT 198.69 65.25 198.89 505.18 ;
      RECT 198.69 65.25 199.29 65.45 ;
      RECT 199.09 63.99 199.29 65.45 ;
      RECT 198.29 65.25 198.49 505.18 ;
      RECT 197.89 65.25 198.49 65.45 ;
      RECT 197.89 63.99 198.09 65.45 ;
      RECT 198.01 58.57 198.21 59.17 ;
      RECT 196.69 58.57 196.89 59.17 ;
      RECT 196.69 58.57 198.21 58.77 ;
      RECT 197.89 37.91 198.09 38.61 ;
      RECT 197.69 37.91 198.09 38.11 ;
      RECT 196.29 63.99 196.49 505.18 ;
      RECT 197.09 63.99 197.29 65.05 ;
      RECT 196.29 63.99 197.29 64.19 ;
      RECT 197.09 65.25 197.29 505.18 ;
      RECT 196.69 65.25 197.29 65.45 ;
      RECT 196.69 64.39 196.89 65.45 ;
      RECT 195.19 510.34 197.19 510.94 ;
      RECT 196.69 65.96 196.89 510.94 ;
      RECT 196.69 37.91 196.89 38.61 ;
      RECT 196.69 37.91 197.09 38.11 ;
      RECT 195.89 63.99 196.09 505.18 ;
      RECT 195.09 63.99 195.29 65.05 ;
      RECT 195.09 63.99 196.09 64.19 ;
      RECT 195.49 37.91 195.69 38.61 ;
      RECT 195.29 37.91 195.69 38.11 ;
      RECT 195.49 58.57 195.69 59.17 ;
      RECT 194.17 58.57 194.37 59.17 ;
      RECT 194.17 58.57 195.69 58.77 ;
      RECT 195.09 65.25 195.29 505.18 ;
      RECT 195.09 65.25 195.69 65.45 ;
      RECT 195.49 64.39 195.69 65.45 ;
      RECT 193.99 510.34 194.79 510.94 ;
      RECT 192.79 510.34 193.59 510.94 ;
      RECT 191.59 510.34 192.39 510.94 ;
      RECT 191.59 510.34 194.79 510.74 ;
      RECT 193.49 68.02 193.69 510.74 ;
      RECT 192.69 68.02 192.89 510.74 ;
      RECT 191.89 65.96 192.09 510.94 ;
      RECT 194.29 37.91 194.49 38.61 ;
      RECT 194.29 37.91 194.69 38.11 ;
      RECT 193.89 65.25 194.09 505.18 ;
      RECT 193.89 65.25 194.49 65.45 ;
      RECT 194.29 63.99 194.49 65.45 ;
      RECT 192.29 65.25 192.49 505.18 ;
      RECT 191.89 65.25 192.49 65.45 ;
      RECT 191.89 63.99 192.09 65.45 ;
      RECT 192.01 58.57 192.21 59.17 ;
      RECT 190.69 58.57 190.89 59.17 ;
      RECT 190.69 58.57 192.21 58.77 ;
      RECT 191.89 37.91 192.09 38.61 ;
      RECT 191.69 37.91 192.09 38.11 ;
      RECT 172.79 38.81 191.49 39.01 ;
      RECT 191.29 37.61 191.49 39.01 ;
      RECT 188.89 37.61 189.09 39.01 ;
      RECT 186.49 37.61 186.69 39.01 ;
      RECT 184.09 37.61 184.29 39.01 ;
      RECT 181.69 37.61 181.89 39.01 ;
      RECT 179.29 37.61 179.49 39.01 ;
      RECT 176.89 37.61 177.09 39.01 ;
      RECT 174.49 37.61 174.69 39.01 ;
      RECT 190.29 63.99 190.49 505.18 ;
      RECT 191.09 63.99 191.29 65.05 ;
      RECT 190.29 63.99 191.29 64.19 ;
      RECT 191.09 65.25 191.29 505.18 ;
      RECT 190.69 65.25 191.29 65.45 ;
      RECT 190.69 64.39 190.89 65.45 ;
      RECT 189.19 510.34 191.19 510.94 ;
      RECT 190.69 65.96 190.89 510.94 ;
      RECT 190.69 37.91 190.89 38.61 ;
      RECT 190.69 37.91 191.09 38.11 ;
      RECT 189.89 63.99 190.09 505.18 ;
      RECT 189.09 63.99 189.29 65.05 ;
      RECT 189.09 63.99 190.09 64.19 ;
      RECT 189.49 37.91 189.69 38.61 ;
      RECT 189.29 37.91 189.69 38.11 ;
      RECT 189.49 58.57 189.69 59.17 ;
      RECT 188.17 58.57 188.37 59.17 ;
      RECT 188.17 58.57 189.69 58.77 ;
      RECT 189.09 65.25 189.29 505.18 ;
      RECT 189.09 65.25 189.69 65.45 ;
      RECT 189.49 64.39 189.69 65.45 ;
      RECT 187.99 510.34 188.79 510.94 ;
      RECT 186.79 510.34 187.59 510.94 ;
      RECT 186.79 510.34 188.79 510.74 ;
      RECT 187.09 65.96 187.29 510.94 ;
      RECT 188.29 37.91 188.49 38.61 ;
      RECT 188.29 37.91 188.69 38.11 ;
      RECT 187.89 65.25 188.09 505.18 ;
      RECT 187.89 65.25 188.49 65.45 ;
      RECT 188.29 63.99 188.49 65.45 ;
      RECT 187.49 65.25 187.69 505.18 ;
      RECT 187.09 65.25 187.69 65.45 ;
      RECT 187.09 63.99 187.29 65.45 ;
      RECT 187.21 58.57 187.41 59.17 ;
      RECT 185.89 58.57 186.09 59.17 ;
      RECT 185.89 58.57 187.41 58.77 ;
      RECT 187.09 37.91 187.29 38.61 ;
      RECT 186.89 37.91 187.29 38.11 ;
      RECT 185.49 63.99 185.69 505.18 ;
      RECT 186.29 63.99 186.49 65.05 ;
      RECT 185.49 63.99 186.49 64.19 ;
      RECT 186.29 65.25 186.49 505.18 ;
      RECT 185.89 65.25 186.49 65.45 ;
      RECT 185.89 64.39 186.09 65.45 ;
      RECT 184.39 510.34 186.39 510.94 ;
      RECT 185.89 65.96 186.09 510.94 ;
      RECT 185.89 37.91 186.09 38.61 ;
      RECT 185.89 37.91 186.29 38.11 ;
      RECT 185.09 63.99 185.29 505.18 ;
      RECT 184.29 63.99 184.49 65.05 ;
      RECT 184.29 63.99 185.29 64.19 ;
      RECT 184.69 37.91 184.89 38.61 ;
      RECT 184.49 37.91 184.89 38.11 ;
      RECT 184.69 58.57 184.89 59.17 ;
      RECT 183.37 58.57 183.57 59.17 ;
      RECT 183.37 58.57 184.89 58.77 ;
      RECT 184.29 65.25 184.49 505.18 ;
      RECT 184.29 65.25 184.89 65.45 ;
      RECT 184.69 64.39 184.89 65.45 ;
      RECT 183.19 510.34 183.99 510.94 ;
      RECT 181.99 510.34 182.79 510.94 ;
      RECT 181.99 510.34 183.99 510.74 ;
      RECT 182.29 65.96 182.49 510.94 ;
      RECT 183.49 37.91 183.69 38.61 ;
      RECT 183.49 37.91 183.89 38.11 ;
      RECT 183.09 65.25 183.29 505.18 ;
      RECT 183.09 65.25 183.69 65.45 ;
      RECT 183.49 63.99 183.69 65.45 ;
      RECT 182.69 65.25 182.89 505.18 ;
      RECT 182.29 65.25 182.89 65.45 ;
      RECT 182.29 63.99 182.49 65.45 ;
      RECT 182.41 58.57 182.61 59.17 ;
      RECT 181.09 58.57 181.29 59.17 ;
      RECT 181.09 58.57 182.61 58.77 ;
      RECT 180.53 24.85 182.59 25.05 ;
      RECT 182.39 24.22 182.59 25.05 ;
      RECT 175.71 12.98 179.39 13.18 ;
      RECT 179.19 12.58 179.39 13.18 ;
      RECT 179.19 12.58 182.49 12.78 ;
      RECT 182.29 37.91 182.49 38.61 ;
      RECT 182.09 37.91 182.49 38.11 ;
      RECT 180.07 23.59 182.45 23.79 ;
      RECT 182.25 22.77 182.45 23.79 ;
      RECT 178.09 22.71 178.29 26.71 ;
      RECT 174.51 22.71 181.87 22.91 ;
      RECT 180.69 63.99 180.89 505.18 ;
      RECT 181.49 63.99 181.69 65.05 ;
      RECT 180.69 63.99 181.69 64.19 ;
      RECT 181.49 65.25 181.69 505.18 ;
      RECT 181.09 65.25 181.69 65.45 ;
      RECT 181.09 64.39 181.29 65.45 ;
      RECT 179.59 510.34 181.59 510.94 ;
      RECT 181.09 65.96 181.29 510.94 ;
      RECT 181.09 37.91 181.29 38.61 ;
      RECT 181.09 37.91 181.49 38.11 ;
      RECT 180.29 63.99 180.49 505.18 ;
      RECT 179.49 63.99 179.69 65.05 ;
      RECT 179.49 63.99 180.49 64.19 ;
      RECT 174.89 16.9 180.46 17.1 ;
      RECT 179.78 15.79 179.98 17.1 ;
      RECT 179.23 15.79 179.98 15.99 ;
      RECT 179.89 37.91 180.09 38.61 ;
      RECT 179.69 37.91 180.09 38.11 ;
      RECT 179.89 58.57 180.09 59.17 ;
      RECT 178.57 58.57 178.77 59.17 ;
      RECT 178.57 58.57 180.09 58.77 ;
      RECT 179.49 65.25 179.69 505.18 ;
      RECT 179.49 65.25 180.09 65.45 ;
      RECT 179.89 64.39 180.09 65.45 ;
      RECT 177.85 16.27 179.58 16.47 ;
      RECT 174.43 16.1 178.05 16.3 ;
      RECT 178.49 23.11 178.69 26.31 ;
      RECT 178.49 23.11 179.29 23.31 ;
      RECT 178.89 26.46 179.29 26.66 ;
      RECT 178.89 24.68 179.09 26.66 ;
      RECT 178.39 510.34 179.19 510.94 ;
      RECT 177.19 510.34 177.99 510.94 ;
      RECT 177.19 510.34 179.19 510.74 ;
      RECT 177.49 65.96 177.69 510.94 ;
      RECT 178.69 37.91 178.89 38.61 ;
      RECT 178.69 37.91 179.09 38.11 ;
      RECT 178.29 65.25 178.49 505.18 ;
      RECT 178.29 65.25 178.89 65.45 ;
      RECT 178.69 63.99 178.89 65.45 ;
      RECT 177.89 65.25 178.09 505.18 ;
      RECT 177.49 65.25 178.09 65.45 ;
      RECT 177.49 63.99 177.69 65.45 ;
      RECT 177.69 23.11 177.89 26.31 ;
      RECT 177.09 23.11 177.89 23.31 ;
      RECT 177.61 58.57 177.81 59.17 ;
      RECT 176.29 58.57 176.49 59.17 ;
      RECT 176.29 58.57 177.81 58.77 ;
      RECT 177.49 37.91 177.69 38.61 ;
      RECT 177.29 37.91 177.69 38.11 ;
      RECT 177.09 26.46 177.49 26.66 ;
      RECT 177.29 24.68 177.49 26.66 ;
      RECT 175.89 63.99 176.09 505.18 ;
      RECT 176.69 63.99 176.89 65.05 ;
      RECT 175.89 63.99 176.89 64.19 ;
      RECT 176.69 65.25 176.89 505.18 ;
      RECT 176.29 65.25 176.89 65.45 ;
      RECT 176.29 64.39 176.49 65.45 ;
      RECT 174.79 510.34 176.79 510.94 ;
      RECT 176.29 65.96 176.49 510.94 ;
      RECT 176.29 37.91 176.49 38.61 ;
      RECT 176.29 37.91 176.69 38.11 ;
      RECT 173.93 23.59 176.31 23.79 ;
      RECT 173.93 22.77 174.13 23.79 ;
      RECT 173.79 24.85 175.85 25.05 ;
      RECT 173.79 24.22 173.99 25.05 ;
      RECT 175.49 63.99 175.69 505.18 ;
      RECT 174.69 63.99 174.89 65.05 ;
      RECT 174.69 63.99 175.69 64.19 ;
      RECT 175.39 15.38 175.59 15.9 ;
      RECT 174.89 15.38 175.59 15.58 ;
      RECT 175.09 37.91 175.29 38.61 ;
      RECT 174.89 37.91 175.29 38.11 ;
      RECT 175.09 58.57 175.29 59.17 ;
      RECT 173.77 58.57 173.97 59.17 ;
      RECT 173.77 58.57 175.29 58.77 ;
      RECT 174.69 65.25 174.89 505.18 ;
      RECT 174.69 65.25 175.29 65.45 ;
      RECT 175.09 64.39 175.29 65.45 ;
      RECT 173.59 510.34 174.39 510.94 ;
      RECT 172.39 510.34 173.19 510.94 ;
      RECT 172.39 510.34 174.39 510.74 ;
      RECT 172.69 65.96 172.89 510.94 ;
      RECT 173.89 37.91 174.09 38.61 ;
      RECT 173.89 37.91 174.29 38.11 ;
      RECT 173.49 65.25 173.69 505.18 ;
      RECT 173.49 65.25 174.09 65.45 ;
      RECT 173.89 63.99 174.09 65.45 ;
      RECT 173.09 65.25 173.29 505.18 ;
      RECT 172.69 65.25 173.29 65.45 ;
      RECT 172.69 63.99 172.89 65.45 ;
      RECT 172.81 58.57 173.01 59.17 ;
      RECT 171.49 58.57 171.69 59.17 ;
      RECT 171.49 58.57 173.01 58.77 ;
      RECT 170.93 24.85 172.99 25.05 ;
      RECT 172.79 24.22 172.99 25.05 ;
      RECT 172.69 37.91 172.89 38.61 ;
      RECT 172.49 37.91 172.89 38.11 ;
      RECT 170.47 23.59 172.85 23.79 ;
      RECT 172.65 22.77 172.85 23.79 ;
      RECT 167.2 16.27 168.93 16.47 ;
      RECT 168.73 16.1 172.35 16.3 ;
      RECT 154.19 38.81 172.29 39.01 ;
      RECT 172.09 37.61 172.29 39.01 ;
      RECT 169.69 37.61 169.89 39.01 ;
      RECT 167.29 37.61 167.49 39.01 ;
      RECT 164.89 37.61 165.09 39.01 ;
      RECT 162.49 37.61 162.69 39.01 ;
      RECT 160.09 37.61 160.29 39.01 ;
      RECT 157.69 37.61 157.89 39.01 ;
      RECT 155.29 37.61 155.49 39.01 ;
      RECT 168.49 22.71 168.69 26.71 ;
      RECT 164.91 22.71 172.27 22.91 ;
      RECT 171.09 63.99 171.29 505.18 ;
      RECT 171.89 63.99 172.09 65.05 ;
      RECT 171.09 63.99 172.09 64.19 ;
      RECT 171.89 65.25 172.09 505.18 ;
      RECT 171.49 65.25 172.09 65.45 ;
      RECT 171.49 64.39 171.69 65.45 ;
      RECT 169.99 510.34 171.99 510.94 ;
      RECT 171.49 65.96 171.69 510.94 ;
      RECT 171.19 15.38 171.39 15.9 ;
      RECT 171.19 15.38 171.89 15.58 ;
      RECT 166.32 16.9 171.89 17.1 ;
      RECT 166.8 15.79 167 17.1 ;
      RECT 166.8 15.79 167.55 15.99 ;
      RECT 171.49 37.91 171.69 38.61 ;
      RECT 171.49 37.91 171.89 38.11 ;
      RECT 167.39 12.98 171.07 13.18 ;
      RECT 167.39 12.58 167.59 13.18 ;
      RECT 164.29 12.58 167.59 12.78 ;
      RECT 170.69 63.99 170.89 505.18 ;
      RECT 169.89 63.99 170.09 65.05 ;
      RECT 169.89 63.99 170.89 64.19 ;
      RECT 170.29 37.91 170.49 38.61 ;
      RECT 170.09 37.91 170.49 38.11 ;
      RECT 170.29 58.57 170.49 59.17 ;
      RECT 168.97 58.57 169.17 59.17 ;
      RECT 168.97 58.57 170.49 58.77 ;
      RECT 169.89 65.25 170.09 505.18 ;
      RECT 169.89 65.25 170.49 65.45 ;
      RECT 170.29 64.39 170.49 65.45 ;
      RECT 168.89 23.11 169.09 26.31 ;
      RECT 168.89 23.11 169.69 23.31 ;
      RECT 169.29 26.46 169.69 26.66 ;
      RECT 169.29 24.68 169.49 26.66 ;
      RECT 168.79 510.34 169.59 510.94 ;
      RECT 167.59 510.34 168.39 510.94 ;
      RECT 167.59 510.34 169.59 510.74 ;
      RECT 167.89 65.96 168.09 510.94 ;
      RECT 169.09 37.91 169.29 38.61 ;
      RECT 169.09 37.91 169.49 38.11 ;
      RECT 168.69 65.25 168.89 505.18 ;
      RECT 168.69 65.25 169.29 65.45 ;
      RECT 169.09 63.99 169.29 65.45 ;
      RECT 168.29 65.25 168.49 505.18 ;
      RECT 167.89 65.25 168.49 65.45 ;
      RECT 167.89 63.99 168.09 65.45 ;
      RECT 168.09 23.11 168.29 26.31 ;
      RECT 167.49 23.11 168.29 23.31 ;
      RECT 168.01 58.57 168.21 59.17 ;
      RECT 166.69 58.57 166.89 59.17 ;
      RECT 166.69 58.57 168.21 58.77 ;
      RECT 167.89 37.91 168.09 38.61 ;
      RECT 167.69 37.91 168.09 38.11 ;
      RECT 167.49 26.46 167.89 26.66 ;
      RECT 167.69 24.68 167.89 26.66 ;
      RECT 166.29 63.99 166.49 505.18 ;
      RECT 167.09 63.99 167.29 65.05 ;
      RECT 166.29 63.99 167.29 64.19 ;
      RECT 167.09 65.25 167.29 505.18 ;
      RECT 166.69 65.25 167.29 65.45 ;
      RECT 166.69 64.39 166.89 65.45 ;
      RECT 165.19 510.34 167.19 510.94 ;
      RECT 166.69 65.96 166.89 510.94 ;
      RECT 166.69 37.91 166.89 38.61 ;
      RECT 166.69 37.91 167.09 38.11 ;
      RECT 164.33 23.59 166.71 23.79 ;
      RECT 164.33 22.77 164.53 23.79 ;
      RECT 164.19 24.85 166.25 25.05 ;
      RECT 164.19 24.22 164.39 25.05 ;
      RECT 165.89 63.99 166.09 505.18 ;
      RECT 165.09 63.99 165.29 65.05 ;
      RECT 165.09 63.99 166.09 64.19 ;
      RECT 165.49 37.91 165.69 38.61 ;
      RECT 165.29 37.91 165.69 38.11 ;
      RECT 165.49 58.57 165.69 59.17 ;
      RECT 164.17 58.57 164.37 59.17 ;
      RECT 164.17 58.57 165.69 58.77 ;
      RECT 165.09 65.25 165.29 505.18 ;
      RECT 165.09 65.25 165.69 65.45 ;
      RECT 165.49 64.39 165.69 65.45 ;
      RECT 163.99 510.34 164.79 510.94 ;
      RECT 162.79 510.34 163.59 510.94 ;
      RECT 162.79 510.34 164.79 510.74 ;
      RECT 163.09 65.96 163.29 510.94 ;
      RECT 164.29 37.91 164.49 38.61 ;
      RECT 164.29 37.91 164.69 38.11 ;
      RECT 163.89 65.25 164.09 505.18 ;
      RECT 163.89 65.25 164.49 65.45 ;
      RECT 164.29 63.99 164.49 65.45 ;
      RECT 163.49 65.25 163.69 505.18 ;
      RECT 163.09 65.25 163.69 65.45 ;
      RECT 163.09 63.99 163.29 65.45 ;
      RECT 163.21 58.57 163.41 59.17 ;
      RECT 161.89 58.57 162.09 59.17 ;
      RECT 161.89 58.57 163.41 58.77 ;
      RECT 163.09 37.91 163.29 38.61 ;
      RECT 162.89 37.91 163.29 38.11 ;
      RECT 161.49 63.99 161.69 505.18 ;
      RECT 162.29 63.99 162.49 65.05 ;
      RECT 161.49 63.99 162.49 64.19 ;
      RECT 162.29 65.25 162.49 505.18 ;
      RECT 161.89 65.25 162.49 65.45 ;
      RECT 161.89 64.39 162.09 65.45 ;
      RECT 160.39 510.34 162.39 510.94 ;
      RECT 161.89 65.96 162.09 510.94 ;
      RECT 161.89 37.91 162.09 38.61 ;
      RECT 161.89 37.91 162.29 38.11 ;
      RECT 161.09 63.99 161.29 505.18 ;
      RECT 160.29 63.99 160.49 65.05 ;
      RECT 160.29 63.99 161.29 64.19 ;
      RECT 160.69 37.91 160.89 38.61 ;
      RECT 160.49 37.91 160.89 38.11 ;
      RECT 160.69 58.57 160.89 59.17 ;
      RECT 159.37 58.57 159.57 59.17 ;
      RECT 159.37 58.57 160.89 58.77 ;
      RECT 160.29 65.25 160.49 505.18 ;
      RECT 160.29 65.25 160.89 65.45 ;
      RECT 160.69 64.39 160.89 65.45 ;
      RECT 159.19 510.34 159.99 510.94 ;
      RECT 157.99 510.34 158.79 510.94 ;
      RECT 157.99 510.34 159.99 510.74 ;
      RECT 158.29 65.96 158.49 510.94 ;
      RECT 159.49 37.91 159.69 38.61 ;
      RECT 159.49 37.91 159.89 38.11 ;
      RECT 159.09 65.25 159.29 505.18 ;
      RECT 159.09 65.25 159.69 65.45 ;
      RECT 159.49 63.99 159.69 65.45 ;
      RECT 158.69 65.25 158.89 505.18 ;
      RECT 158.29 65.25 158.89 65.45 ;
      RECT 158.29 63.99 158.49 65.45 ;
      RECT 158.41 58.57 158.61 59.17 ;
      RECT 157.09 58.57 157.29 59.17 ;
      RECT 157.09 58.57 158.61 58.77 ;
      RECT 158.29 37.91 158.49 38.61 ;
      RECT 158.09 37.91 158.49 38.11 ;
      RECT 156.69 63.99 156.89 505.18 ;
      RECT 157.49 63.99 157.69 65.05 ;
      RECT 156.69 63.99 157.69 64.19 ;
      RECT 157.49 65.25 157.69 505.18 ;
      RECT 157.09 65.25 157.69 65.45 ;
      RECT 157.09 64.39 157.29 65.45 ;
      RECT 155.59 510.34 157.59 510.94 ;
      RECT 157.09 65.96 157.29 510.94 ;
      RECT 157.09 37.91 157.29 38.61 ;
      RECT 157.09 37.91 157.49 38.11 ;
      RECT 156.29 63.99 156.49 505.18 ;
      RECT 155.49 63.99 155.69 65.05 ;
      RECT 155.49 63.99 156.49 64.19 ;
      RECT 155.89 37.91 156.09 38.61 ;
      RECT 155.69 37.91 156.09 38.11 ;
      RECT 155.89 58.57 156.09 59.17 ;
      RECT 154.57 58.57 154.77 59.17 ;
      RECT 154.57 58.57 156.09 58.77 ;
      RECT 155.49 65.25 155.69 505.18 ;
      RECT 155.49 65.25 156.09 65.45 ;
      RECT 155.89 64.39 156.09 65.45 ;
      RECT 154.39 510.34 155.19 510.94 ;
      RECT 153.19 510.34 153.99 510.94 ;
      RECT 153.19 510.34 155.19 510.74 ;
      RECT 153.09 67.66 153.29 510.54 ;
      RECT 153.89 67.66 154.09 510.74 ;
      RECT 153.09 67.66 154.09 67.86 ;
      RECT 154.69 37.91 154.89 38.61 ;
      RECT 154.69 37.91 155.09 38.11 ;
      RECT 154.29 65.25 154.49 505.18 ;
      RECT 154.29 65.25 154.89 65.45 ;
      RECT 154.69 63.99 154.89 65.45 ;
      RECT 142.6 30.35 153.09 30.55 ;
      RECT 147.69 30.21 148.04 30.55 ;
      RECT 123.2 66.83 126.04 68.11 ;
      RECT 123.2 66.83 152.69 67.63 ;
      RECT 149.11 65.83 150.15 67.63 ;
      RECT 147.19 65.83 148.23 67.63 ;
      RECT 145.27 65.83 146.31 67.63 ;
      RECT 143.35 65.83 144.39 67.63 ;
      RECT 86.81 28.01 141.59 30.21 ;
      RECT 86.81 28.31 151.37 29.15 ;
      RECT 86.81 28.01 144.77 29.15 ;
      RECT 150.21 507.13 150.41 509 ;
      RECT 149.71 507.13 150.41 507.33 ;
      RECT 149.71 506.34 149.93 507.33 ;
      RECT 114.94 506.74 137.41 506.94 ;
      RECT 137.21 506.34 137.41 506.94 ;
      RECT 137.21 506.34 149.93 506.54 ;
      RECT 147.95 69.86 148.55 71.1 ;
      RECT 147.95 70.16 150.33 70.66 ;
      RECT 109.46 69.86 148.55 70.16 ;
      RECT 109.46 72.36 148.55 72.66 ;
      RECT 147.95 71.42 148.55 72.66 ;
      RECT 147.95 71.86 150.33 72.36 ;
      RECT 147.95 73.26 148.55 74.5 ;
      RECT 147.95 73.56 150.33 74.06 ;
      RECT 109.46 73.26 148.55 73.56 ;
      RECT 109.46 75.76 148.55 76.06 ;
      RECT 147.95 74.82 148.55 76.06 ;
      RECT 147.95 75.26 150.33 75.76 ;
      RECT 147.95 76.66 148.55 77.9 ;
      RECT 147.95 76.96 150.33 77.46 ;
      RECT 109.46 76.66 148.55 76.96 ;
      RECT 109.46 79.16 148.55 79.46 ;
      RECT 147.95 78.22 148.55 79.46 ;
      RECT 147.95 78.66 150.33 79.16 ;
      RECT 147.95 80.06 148.55 81.3 ;
      RECT 147.95 80.36 150.33 80.86 ;
      RECT 109.46 80.06 148.55 80.36 ;
      RECT 109.46 82.56 148.55 82.86 ;
      RECT 147.95 81.62 148.55 82.86 ;
      RECT 147.95 82.06 150.33 82.56 ;
      RECT 147.95 83.46 148.55 84.7 ;
      RECT 147.95 83.76 150.33 84.26 ;
      RECT 109.46 83.46 148.55 83.76 ;
      RECT 109.46 85.96 148.55 86.26 ;
      RECT 147.95 85.02 148.55 86.26 ;
      RECT 147.95 85.46 150.33 85.96 ;
      RECT 147.95 86.86 148.55 88.1 ;
      RECT 147.95 87.16 150.33 87.66 ;
      RECT 109.46 86.86 148.55 87.16 ;
      RECT 109.46 89.36 148.55 89.66 ;
      RECT 147.95 88.42 148.55 89.66 ;
      RECT 147.95 88.86 150.33 89.36 ;
      RECT 147.95 90.26 148.55 91.5 ;
      RECT 147.95 90.56 150.33 91.06 ;
      RECT 109.46 90.26 148.55 90.56 ;
      RECT 109.46 92.76 148.55 93.06 ;
      RECT 147.95 91.82 148.55 93.06 ;
      RECT 147.95 92.26 150.33 92.76 ;
      RECT 147.95 93.66 148.55 94.9 ;
      RECT 147.95 93.96 150.33 94.46 ;
      RECT 109.46 93.66 148.55 93.96 ;
      RECT 109.46 96.16 148.55 96.46 ;
      RECT 147.95 95.22 148.55 96.46 ;
      RECT 147.95 95.66 150.33 96.16 ;
      RECT 147.95 97.06 148.55 98.3 ;
      RECT 147.95 97.36 150.33 97.86 ;
      RECT 109.46 97.06 148.55 97.36 ;
      RECT 109.46 99.56 148.55 99.86 ;
      RECT 147.95 98.62 148.55 99.86 ;
      RECT 147.95 99.06 150.33 99.56 ;
      RECT 147.95 100.46 148.55 101.7 ;
      RECT 147.95 100.76 150.33 101.26 ;
      RECT 109.46 100.46 148.55 100.76 ;
      RECT 109.46 102.96 148.55 103.26 ;
      RECT 147.95 102.02 148.55 103.26 ;
      RECT 147.95 102.46 150.33 102.96 ;
      RECT 147.95 103.86 148.55 105.1 ;
      RECT 147.95 104.16 150.33 104.66 ;
      RECT 109.46 103.86 148.55 104.16 ;
      RECT 109.46 106.36 148.55 106.66 ;
      RECT 147.95 105.42 148.55 106.66 ;
      RECT 147.95 105.86 150.33 106.36 ;
      RECT 147.95 107.26 148.55 108.5 ;
      RECT 147.95 107.56 150.33 108.06 ;
      RECT 109.46 107.26 148.55 107.56 ;
      RECT 109.46 109.76 148.55 110.06 ;
      RECT 147.95 108.82 148.55 110.06 ;
      RECT 147.95 109.26 150.33 109.76 ;
      RECT 147.95 110.66 148.55 111.9 ;
      RECT 147.95 110.96 150.33 111.46 ;
      RECT 109.46 110.66 148.55 110.96 ;
      RECT 109.46 113.16 148.55 113.46 ;
      RECT 147.95 112.22 148.55 113.46 ;
      RECT 147.95 112.66 150.33 113.16 ;
      RECT 147.95 114.06 148.55 115.3 ;
      RECT 147.95 114.36 150.33 114.86 ;
      RECT 109.46 114.06 148.55 114.36 ;
      RECT 109.46 116.56 148.55 116.86 ;
      RECT 147.95 115.62 148.55 116.86 ;
      RECT 147.95 116.06 150.33 116.56 ;
      RECT 147.95 117.46 148.55 118.7 ;
      RECT 147.95 117.76 150.33 118.26 ;
      RECT 109.46 117.46 148.55 117.76 ;
      RECT 109.46 119.96 148.55 120.26 ;
      RECT 147.95 119.02 148.55 120.26 ;
      RECT 147.95 119.46 150.33 119.96 ;
      RECT 147.95 120.86 148.55 122.1 ;
      RECT 147.95 121.16 150.33 121.66 ;
      RECT 109.46 120.86 148.55 121.16 ;
      RECT 109.46 123.36 148.55 123.66 ;
      RECT 147.95 122.42 148.55 123.66 ;
      RECT 147.95 122.86 150.33 123.36 ;
      RECT 147.95 124.26 148.55 125.5 ;
      RECT 147.95 124.56 150.33 125.06 ;
      RECT 109.46 124.26 148.55 124.56 ;
      RECT 109.46 126.76 148.55 127.06 ;
      RECT 147.95 125.82 148.55 127.06 ;
      RECT 147.95 126.26 150.33 126.76 ;
      RECT 147.95 127.66 148.55 128.9 ;
      RECT 147.95 127.96 150.33 128.46 ;
      RECT 109.46 127.66 148.55 127.96 ;
      RECT 109.46 130.16 148.55 130.46 ;
      RECT 147.95 129.22 148.55 130.46 ;
      RECT 147.95 129.66 150.33 130.16 ;
      RECT 147.95 131.06 148.55 132.3 ;
      RECT 147.95 131.36 150.33 131.86 ;
      RECT 109.46 131.06 148.55 131.36 ;
      RECT 109.46 133.56 148.55 133.86 ;
      RECT 147.95 132.62 148.55 133.86 ;
      RECT 147.95 133.06 150.33 133.56 ;
      RECT 147.95 134.46 148.55 135.7 ;
      RECT 147.95 134.76 150.33 135.26 ;
      RECT 109.46 134.46 148.55 134.76 ;
      RECT 109.46 136.96 148.55 137.26 ;
      RECT 147.95 136.02 148.55 137.26 ;
      RECT 147.95 136.46 150.33 136.96 ;
      RECT 147.95 137.86 148.55 139.1 ;
      RECT 147.95 138.16 150.33 138.66 ;
      RECT 109.46 137.86 148.55 138.16 ;
      RECT 109.46 140.36 148.55 140.66 ;
      RECT 147.95 139.42 148.55 140.66 ;
      RECT 147.95 139.86 150.33 140.36 ;
      RECT 147.95 141.26 148.55 142.5 ;
      RECT 147.95 141.56 150.33 142.06 ;
      RECT 109.46 141.26 148.55 141.56 ;
      RECT 109.46 143.76 148.55 144.06 ;
      RECT 147.95 142.82 148.55 144.06 ;
      RECT 147.95 143.26 150.33 143.76 ;
      RECT 147.95 144.66 148.55 145.9 ;
      RECT 147.95 144.96 150.33 145.46 ;
      RECT 109.46 144.66 148.55 144.96 ;
      RECT 109.46 147.16 148.55 147.46 ;
      RECT 147.95 146.22 148.55 147.46 ;
      RECT 147.95 146.66 150.33 147.16 ;
      RECT 147.95 148.06 148.55 149.3 ;
      RECT 147.95 148.36 150.33 148.86 ;
      RECT 109.46 148.06 148.55 148.36 ;
      RECT 109.46 150.56 148.55 150.86 ;
      RECT 147.95 149.62 148.55 150.86 ;
      RECT 147.95 150.06 150.33 150.56 ;
      RECT 147.95 151.46 148.55 152.7 ;
      RECT 147.95 151.76 150.33 152.26 ;
      RECT 109.46 151.46 148.55 151.76 ;
      RECT 109.46 153.96 148.55 154.26 ;
      RECT 147.95 153.02 148.55 154.26 ;
      RECT 147.95 153.46 150.33 153.96 ;
      RECT 147.95 154.86 148.55 156.1 ;
      RECT 147.95 155.16 150.33 155.66 ;
      RECT 109.46 154.86 148.55 155.16 ;
      RECT 109.46 157.36 148.55 157.66 ;
      RECT 147.95 156.42 148.55 157.66 ;
      RECT 147.95 156.86 150.33 157.36 ;
      RECT 147.95 158.26 148.55 159.5 ;
      RECT 147.95 158.56 150.33 159.06 ;
      RECT 109.46 158.26 148.55 158.56 ;
      RECT 109.46 160.76 148.55 161.06 ;
      RECT 147.95 159.82 148.55 161.06 ;
      RECT 147.95 160.26 150.33 160.76 ;
      RECT 147.95 161.66 148.55 162.9 ;
      RECT 147.95 161.96 150.33 162.46 ;
      RECT 109.46 161.66 148.55 161.96 ;
      RECT 109.46 164.16 148.55 164.46 ;
      RECT 147.95 163.22 148.55 164.46 ;
      RECT 147.95 163.66 150.33 164.16 ;
      RECT 147.95 165.06 148.55 166.3 ;
      RECT 147.95 165.36 150.33 165.86 ;
      RECT 109.46 165.06 148.55 165.36 ;
      RECT 109.46 167.56 148.55 167.86 ;
      RECT 147.95 166.62 148.55 167.86 ;
      RECT 147.95 167.06 150.33 167.56 ;
      RECT 147.95 168.46 148.55 169.7 ;
      RECT 147.95 168.76 150.33 169.26 ;
      RECT 109.46 168.46 148.55 168.76 ;
      RECT 109.46 170.96 148.55 171.26 ;
      RECT 147.95 170.02 148.55 171.26 ;
      RECT 147.95 170.46 150.33 170.96 ;
      RECT 147.95 171.86 148.55 173.1 ;
      RECT 147.95 172.16 150.33 172.66 ;
      RECT 109.46 171.86 148.55 172.16 ;
      RECT 109.46 174.36 148.55 174.66 ;
      RECT 147.95 173.42 148.55 174.66 ;
      RECT 147.95 173.86 150.33 174.36 ;
      RECT 147.95 175.26 148.55 176.5 ;
      RECT 147.95 175.56 150.33 176.06 ;
      RECT 109.46 175.26 148.55 175.56 ;
      RECT 109.46 177.76 148.55 178.06 ;
      RECT 147.95 176.82 148.55 178.06 ;
      RECT 147.95 177.26 150.33 177.76 ;
      RECT 147.95 178.66 148.55 179.9 ;
      RECT 147.95 178.96 150.33 179.46 ;
      RECT 109.46 178.66 148.55 178.96 ;
      RECT 109.46 181.16 148.55 181.46 ;
      RECT 147.95 180.22 148.55 181.46 ;
      RECT 147.95 180.66 150.33 181.16 ;
      RECT 147.95 182.06 148.55 183.3 ;
      RECT 147.95 182.36 150.33 182.86 ;
      RECT 109.46 182.06 148.55 182.36 ;
      RECT 109.46 184.56 148.55 184.86 ;
      RECT 147.95 183.62 148.55 184.86 ;
      RECT 147.95 184.06 150.33 184.56 ;
      RECT 147.95 185.46 148.55 186.7 ;
      RECT 147.95 185.76 150.33 186.26 ;
      RECT 109.46 185.46 148.55 185.76 ;
      RECT 109.46 187.96 148.55 188.26 ;
      RECT 147.95 187.02 148.55 188.26 ;
      RECT 147.95 187.46 150.33 187.96 ;
      RECT 147.95 188.86 148.55 190.1 ;
      RECT 147.95 189.16 150.33 189.66 ;
      RECT 109.46 188.86 148.55 189.16 ;
      RECT 109.46 191.36 148.55 191.66 ;
      RECT 147.95 190.42 148.55 191.66 ;
      RECT 147.95 190.86 150.33 191.36 ;
      RECT 147.95 192.26 148.55 193.5 ;
      RECT 147.95 192.56 150.33 193.06 ;
      RECT 109.46 192.26 148.55 192.56 ;
      RECT 109.46 194.76 148.55 195.06 ;
      RECT 147.95 193.82 148.55 195.06 ;
      RECT 147.95 194.26 150.33 194.76 ;
      RECT 147.95 195.66 148.55 196.9 ;
      RECT 147.95 195.96 150.33 196.46 ;
      RECT 109.46 195.66 148.55 195.96 ;
      RECT 109.46 198.16 148.55 198.46 ;
      RECT 147.95 197.22 148.55 198.46 ;
      RECT 147.95 197.66 150.33 198.16 ;
      RECT 147.95 199.06 148.55 200.3 ;
      RECT 147.95 199.36 150.33 199.86 ;
      RECT 109.46 199.06 148.55 199.36 ;
      RECT 109.46 201.56 148.55 201.86 ;
      RECT 147.95 200.62 148.55 201.86 ;
      RECT 147.95 201.06 150.33 201.56 ;
      RECT 147.95 202.46 148.55 203.7 ;
      RECT 147.95 202.76 150.33 203.26 ;
      RECT 109.46 202.46 148.55 202.76 ;
      RECT 109.46 204.96 148.55 205.26 ;
      RECT 147.95 204.02 148.55 205.26 ;
      RECT 147.95 204.46 150.33 204.96 ;
      RECT 147.95 205.86 148.55 207.1 ;
      RECT 147.95 206.16 150.33 206.66 ;
      RECT 109.46 205.86 148.55 206.16 ;
      RECT 109.46 208.36 148.55 208.66 ;
      RECT 147.95 207.42 148.55 208.66 ;
      RECT 147.95 207.86 150.33 208.36 ;
      RECT 147.95 209.26 148.55 210.5 ;
      RECT 147.95 209.56 150.33 210.06 ;
      RECT 109.46 209.26 148.55 209.56 ;
      RECT 109.46 211.76 148.55 212.06 ;
      RECT 147.95 210.82 148.55 212.06 ;
      RECT 147.95 211.26 150.33 211.76 ;
      RECT 147.95 212.66 148.55 213.9 ;
      RECT 147.95 212.96 150.33 213.46 ;
      RECT 109.46 212.66 148.55 212.96 ;
      RECT 109.46 215.16 148.55 215.46 ;
      RECT 147.95 214.22 148.55 215.46 ;
      RECT 147.95 214.66 150.33 215.16 ;
      RECT 147.95 216.06 148.55 217.3 ;
      RECT 147.95 216.36 150.33 216.86 ;
      RECT 109.46 216.06 148.55 216.36 ;
      RECT 109.46 218.56 148.55 218.86 ;
      RECT 147.95 217.62 148.55 218.86 ;
      RECT 147.95 218.06 150.33 218.56 ;
      RECT 147.95 219.46 148.55 220.7 ;
      RECT 147.95 219.76 150.33 220.26 ;
      RECT 109.46 219.46 148.55 219.76 ;
      RECT 109.46 221.96 148.55 222.26 ;
      RECT 147.95 221.02 148.55 222.26 ;
      RECT 147.95 221.46 150.33 221.96 ;
      RECT 147.95 222.86 148.55 224.1 ;
      RECT 147.95 223.16 150.33 223.66 ;
      RECT 109.46 222.86 148.55 223.16 ;
      RECT 109.46 225.36 148.55 225.66 ;
      RECT 147.95 224.42 148.55 225.66 ;
      RECT 147.95 224.86 150.33 225.36 ;
      RECT 147.95 226.26 148.55 227.5 ;
      RECT 147.95 226.56 150.33 227.06 ;
      RECT 109.46 226.26 148.55 226.56 ;
      RECT 109.46 228.76 148.55 229.06 ;
      RECT 147.95 227.82 148.55 229.06 ;
      RECT 147.95 228.26 150.33 228.76 ;
      RECT 147.95 229.66 148.55 230.9 ;
      RECT 147.95 229.96 150.33 230.46 ;
      RECT 109.46 229.66 148.55 229.96 ;
      RECT 109.46 232.16 148.55 232.46 ;
      RECT 147.95 231.22 148.55 232.46 ;
      RECT 147.95 231.66 150.33 232.16 ;
      RECT 147.95 233.06 148.55 234.3 ;
      RECT 147.95 233.36 150.33 233.86 ;
      RECT 109.46 233.06 148.55 233.36 ;
      RECT 109.46 235.56 148.55 235.86 ;
      RECT 147.95 234.62 148.55 235.86 ;
      RECT 147.95 235.06 150.33 235.56 ;
      RECT 147.95 236.46 148.55 237.7 ;
      RECT 147.95 236.76 150.33 237.26 ;
      RECT 109.46 236.46 148.55 236.76 ;
      RECT 109.46 238.96 148.55 239.26 ;
      RECT 147.95 238.02 148.55 239.26 ;
      RECT 147.95 238.46 150.33 238.96 ;
      RECT 147.95 239.86 148.55 241.1 ;
      RECT 147.95 240.16 150.33 240.66 ;
      RECT 109.46 239.86 148.55 240.16 ;
      RECT 109.46 242.36 148.55 242.66 ;
      RECT 147.95 241.42 148.55 242.66 ;
      RECT 147.95 241.86 150.33 242.36 ;
      RECT 147.95 243.26 148.55 244.5 ;
      RECT 147.95 243.56 150.33 244.06 ;
      RECT 109.46 243.26 148.55 243.56 ;
      RECT 109.46 245.76 148.55 246.06 ;
      RECT 147.95 244.82 148.55 246.06 ;
      RECT 147.95 245.26 150.33 245.76 ;
      RECT 147.95 246.66 148.55 247.9 ;
      RECT 147.95 246.96 150.33 247.46 ;
      RECT 109.46 246.66 148.55 246.96 ;
      RECT 109.46 249.16 148.55 249.46 ;
      RECT 147.95 248.22 148.55 249.46 ;
      RECT 147.95 248.66 150.33 249.16 ;
      RECT 147.95 250.06 148.55 251.3 ;
      RECT 147.95 250.36 150.33 250.86 ;
      RECT 109.46 250.06 148.55 250.36 ;
      RECT 109.46 252.56 148.55 252.86 ;
      RECT 147.95 251.62 148.55 252.86 ;
      RECT 147.95 252.06 150.33 252.56 ;
      RECT 147.95 253.46 148.55 254.7 ;
      RECT 147.95 253.76 150.33 254.26 ;
      RECT 109.46 253.46 148.55 253.76 ;
      RECT 109.46 255.96 148.55 256.26 ;
      RECT 147.95 255.02 148.55 256.26 ;
      RECT 147.95 255.46 150.33 255.96 ;
      RECT 147.95 256.86 148.55 258.1 ;
      RECT 147.95 257.16 150.33 257.66 ;
      RECT 109.46 256.86 148.55 257.16 ;
      RECT 109.46 259.36 148.55 259.66 ;
      RECT 147.95 258.42 148.55 259.66 ;
      RECT 147.95 258.86 150.33 259.36 ;
      RECT 147.95 260.26 148.55 261.5 ;
      RECT 147.95 260.56 150.33 261.06 ;
      RECT 109.46 260.26 148.55 260.56 ;
      RECT 109.46 262.76 148.55 263.06 ;
      RECT 147.95 261.82 148.55 263.06 ;
      RECT 147.95 262.26 150.33 262.76 ;
      RECT 147.95 263.66 148.55 264.9 ;
      RECT 147.95 263.96 150.33 264.46 ;
      RECT 109.46 263.66 148.55 263.96 ;
      RECT 109.46 266.16 148.55 266.46 ;
      RECT 147.95 265.22 148.55 266.46 ;
      RECT 147.95 265.66 150.33 266.16 ;
      RECT 147.95 267.06 148.55 268.3 ;
      RECT 147.95 267.36 150.33 267.86 ;
      RECT 109.46 267.06 148.55 267.36 ;
      RECT 109.46 269.56 148.55 269.86 ;
      RECT 147.95 268.62 148.55 269.86 ;
      RECT 147.95 269.06 150.33 269.56 ;
      RECT 147.95 270.46 148.55 271.7 ;
      RECT 147.95 270.76 150.33 271.26 ;
      RECT 109.46 270.46 148.55 270.76 ;
      RECT 109.46 272.96 148.55 273.26 ;
      RECT 147.95 272.02 148.55 273.26 ;
      RECT 147.95 272.46 150.33 272.96 ;
      RECT 147.95 273.86 148.55 275.1 ;
      RECT 147.95 274.16 150.33 274.66 ;
      RECT 109.46 273.86 148.55 274.16 ;
      RECT 109.46 276.36 148.55 276.66 ;
      RECT 147.95 275.42 148.55 276.66 ;
      RECT 147.95 275.86 150.33 276.36 ;
      RECT 147.95 277.26 148.55 278.5 ;
      RECT 147.95 277.56 150.33 278.06 ;
      RECT 109.46 277.26 148.55 277.56 ;
      RECT 109.46 279.76 148.55 280.06 ;
      RECT 147.95 278.82 148.55 280.06 ;
      RECT 147.95 279.26 150.33 279.76 ;
      RECT 147.95 280.66 148.55 281.9 ;
      RECT 147.95 280.96 150.33 281.46 ;
      RECT 109.46 280.66 148.55 280.96 ;
      RECT 109.46 283.16 148.55 283.46 ;
      RECT 147.95 282.22 148.55 283.46 ;
      RECT 147.95 282.66 150.33 283.16 ;
      RECT 147.95 284.06 148.55 285.3 ;
      RECT 147.95 284.36 150.33 284.86 ;
      RECT 109.46 284.06 148.55 284.36 ;
      RECT 109.46 286.56 148.55 286.86 ;
      RECT 147.95 285.62 148.55 286.86 ;
      RECT 147.95 286.06 150.33 286.56 ;
      RECT 147.95 287.46 148.55 288.7 ;
      RECT 147.95 287.76 150.33 288.26 ;
      RECT 109.46 287.46 148.55 287.76 ;
      RECT 109.46 289.96 148.55 290.26 ;
      RECT 147.95 289.02 148.55 290.26 ;
      RECT 147.95 289.46 150.33 289.96 ;
      RECT 147.95 290.86 148.55 292.1 ;
      RECT 147.95 291.16 150.33 291.66 ;
      RECT 109.46 290.86 148.55 291.16 ;
      RECT 109.46 293.36 148.55 293.66 ;
      RECT 147.95 292.42 148.55 293.66 ;
      RECT 147.95 292.86 150.33 293.36 ;
      RECT 147.95 294.26 148.55 295.5 ;
      RECT 147.95 294.56 150.33 295.06 ;
      RECT 109.46 294.26 148.55 294.56 ;
      RECT 109.46 296.76 148.55 297.06 ;
      RECT 147.95 295.82 148.55 297.06 ;
      RECT 147.95 296.26 150.33 296.76 ;
      RECT 147.95 297.66 148.55 298.9 ;
      RECT 147.95 297.96 150.33 298.46 ;
      RECT 109.46 297.66 148.55 297.96 ;
      RECT 109.46 300.16 148.55 300.46 ;
      RECT 147.95 299.22 148.55 300.46 ;
      RECT 147.95 299.66 150.33 300.16 ;
      RECT 147.95 301.06 148.55 302.3 ;
      RECT 147.95 301.36 150.33 301.86 ;
      RECT 109.46 301.06 148.55 301.36 ;
      RECT 109.46 303.56 148.55 303.86 ;
      RECT 147.95 302.62 148.55 303.86 ;
      RECT 147.95 303.06 150.33 303.56 ;
      RECT 147.95 304.46 148.55 305.7 ;
      RECT 147.95 304.76 150.33 305.26 ;
      RECT 109.46 304.46 148.55 304.76 ;
      RECT 109.46 306.96 148.55 307.26 ;
      RECT 147.95 306.02 148.55 307.26 ;
      RECT 147.95 306.46 150.33 306.96 ;
      RECT 147.95 307.86 148.55 309.1 ;
      RECT 147.95 308.16 150.33 308.66 ;
      RECT 109.46 307.86 148.55 308.16 ;
      RECT 109.46 310.36 148.55 310.66 ;
      RECT 147.95 309.42 148.55 310.66 ;
      RECT 147.95 309.86 150.33 310.36 ;
      RECT 147.95 311.26 148.55 312.5 ;
      RECT 147.95 311.56 150.33 312.06 ;
      RECT 109.46 311.26 148.55 311.56 ;
      RECT 109.46 313.76 148.55 314.06 ;
      RECT 147.95 312.82 148.55 314.06 ;
      RECT 147.95 313.26 150.33 313.76 ;
      RECT 147.95 314.66 148.55 315.9 ;
      RECT 147.95 314.96 150.33 315.46 ;
      RECT 109.46 314.66 148.55 314.96 ;
      RECT 109.46 317.16 148.55 317.46 ;
      RECT 147.95 316.22 148.55 317.46 ;
      RECT 147.95 316.66 150.33 317.16 ;
      RECT 147.95 318.06 148.55 319.3 ;
      RECT 147.95 318.36 150.33 318.86 ;
      RECT 109.46 318.06 148.55 318.36 ;
      RECT 109.46 320.56 148.55 320.86 ;
      RECT 147.95 319.62 148.55 320.86 ;
      RECT 147.95 320.06 150.33 320.56 ;
      RECT 147.95 321.46 148.55 322.7 ;
      RECT 147.95 321.76 150.33 322.26 ;
      RECT 109.46 321.46 148.55 321.76 ;
      RECT 109.46 323.96 148.55 324.26 ;
      RECT 147.95 323.02 148.55 324.26 ;
      RECT 147.95 323.46 150.33 323.96 ;
      RECT 147.95 324.86 148.55 326.1 ;
      RECT 147.95 325.16 150.33 325.66 ;
      RECT 109.46 324.86 148.55 325.16 ;
      RECT 109.46 327.36 148.55 327.66 ;
      RECT 147.95 326.42 148.55 327.66 ;
      RECT 147.95 326.86 150.33 327.36 ;
      RECT 147.95 328.26 148.55 329.5 ;
      RECT 147.95 328.56 150.33 329.06 ;
      RECT 109.46 328.26 148.55 328.56 ;
      RECT 109.46 330.76 148.55 331.06 ;
      RECT 147.95 329.82 148.55 331.06 ;
      RECT 147.95 330.26 150.33 330.76 ;
      RECT 147.95 331.66 148.55 332.9 ;
      RECT 147.95 331.96 150.33 332.46 ;
      RECT 109.46 331.66 148.55 331.96 ;
      RECT 109.46 334.16 148.55 334.46 ;
      RECT 147.95 333.22 148.55 334.46 ;
      RECT 147.95 333.66 150.33 334.16 ;
      RECT 147.95 335.06 148.55 336.3 ;
      RECT 147.95 335.36 150.33 335.86 ;
      RECT 109.46 335.06 148.55 335.36 ;
      RECT 109.46 337.56 148.55 337.86 ;
      RECT 147.95 336.62 148.55 337.86 ;
      RECT 147.95 337.06 150.33 337.56 ;
      RECT 147.95 338.46 148.55 339.7 ;
      RECT 147.95 338.76 150.33 339.26 ;
      RECT 109.46 338.46 148.55 338.76 ;
      RECT 109.46 340.96 148.55 341.26 ;
      RECT 147.95 340.02 148.55 341.26 ;
      RECT 147.95 340.46 150.33 340.96 ;
      RECT 147.95 341.86 148.55 343.1 ;
      RECT 147.95 342.16 150.33 342.66 ;
      RECT 109.46 341.86 148.55 342.16 ;
      RECT 109.46 344.36 148.55 344.66 ;
      RECT 147.95 343.42 148.55 344.66 ;
      RECT 147.95 343.86 150.33 344.36 ;
      RECT 147.95 345.26 148.55 346.5 ;
      RECT 147.95 345.56 150.33 346.06 ;
      RECT 109.46 345.26 148.55 345.56 ;
      RECT 109.46 347.76 148.55 348.06 ;
      RECT 147.95 346.82 148.55 348.06 ;
      RECT 147.95 347.26 150.33 347.76 ;
      RECT 147.95 348.66 148.55 349.9 ;
      RECT 147.95 348.96 150.33 349.46 ;
      RECT 109.46 348.66 148.55 348.96 ;
      RECT 109.46 351.16 148.55 351.46 ;
      RECT 147.95 350.22 148.55 351.46 ;
      RECT 147.95 350.66 150.33 351.16 ;
      RECT 147.95 352.06 148.55 353.3 ;
      RECT 147.95 352.36 150.33 352.86 ;
      RECT 109.46 352.06 148.55 352.36 ;
      RECT 109.46 354.56 148.55 354.86 ;
      RECT 147.95 353.62 148.55 354.86 ;
      RECT 147.95 354.06 150.33 354.56 ;
      RECT 147.95 355.46 148.55 356.7 ;
      RECT 147.95 355.76 150.33 356.26 ;
      RECT 109.46 355.46 148.55 355.76 ;
      RECT 109.46 357.96 148.55 358.26 ;
      RECT 147.95 357.02 148.55 358.26 ;
      RECT 147.95 357.46 150.33 357.96 ;
      RECT 147.95 358.86 148.55 360.1 ;
      RECT 147.95 359.16 150.33 359.66 ;
      RECT 109.46 358.86 148.55 359.16 ;
      RECT 109.46 361.36 148.55 361.66 ;
      RECT 147.95 360.42 148.55 361.66 ;
      RECT 147.95 360.86 150.33 361.36 ;
      RECT 147.95 362.26 148.55 363.5 ;
      RECT 147.95 362.56 150.33 363.06 ;
      RECT 109.46 362.26 148.55 362.56 ;
      RECT 109.46 364.76 148.55 365.06 ;
      RECT 147.95 363.82 148.55 365.06 ;
      RECT 147.95 364.26 150.33 364.76 ;
      RECT 147.95 365.66 148.55 366.9 ;
      RECT 147.95 365.96 150.33 366.46 ;
      RECT 109.46 365.66 148.55 365.96 ;
      RECT 109.46 368.16 148.55 368.46 ;
      RECT 147.95 367.22 148.55 368.46 ;
      RECT 147.95 367.66 150.33 368.16 ;
      RECT 147.95 369.06 148.55 370.3 ;
      RECT 147.95 369.36 150.33 369.86 ;
      RECT 109.46 369.06 148.55 369.36 ;
      RECT 109.46 371.56 148.55 371.86 ;
      RECT 147.95 370.62 148.55 371.86 ;
      RECT 147.95 371.06 150.33 371.56 ;
      RECT 147.95 372.46 148.55 373.7 ;
      RECT 147.95 372.76 150.33 373.26 ;
      RECT 109.46 372.46 148.55 372.76 ;
      RECT 109.46 374.96 148.55 375.26 ;
      RECT 147.95 374.02 148.55 375.26 ;
      RECT 147.95 374.46 150.33 374.96 ;
      RECT 147.95 375.86 148.55 377.1 ;
      RECT 147.95 376.16 150.33 376.66 ;
      RECT 109.46 375.86 148.55 376.16 ;
      RECT 109.46 378.36 148.55 378.66 ;
      RECT 147.95 377.42 148.55 378.66 ;
      RECT 147.95 377.86 150.33 378.36 ;
      RECT 147.95 379.26 148.55 380.5 ;
      RECT 147.95 379.56 150.33 380.06 ;
      RECT 109.46 379.26 148.55 379.56 ;
      RECT 109.46 381.76 148.55 382.06 ;
      RECT 147.95 380.82 148.55 382.06 ;
      RECT 147.95 381.26 150.33 381.76 ;
      RECT 147.95 382.66 148.55 383.9 ;
      RECT 147.95 382.96 150.33 383.46 ;
      RECT 109.46 382.66 148.55 382.96 ;
      RECT 109.46 385.16 148.55 385.46 ;
      RECT 147.95 384.22 148.55 385.46 ;
      RECT 147.95 384.66 150.33 385.16 ;
      RECT 147.95 386.06 148.55 387.3 ;
      RECT 147.95 386.36 150.33 386.86 ;
      RECT 109.46 386.06 148.55 386.36 ;
      RECT 109.46 388.56 148.55 388.86 ;
      RECT 147.95 387.62 148.55 388.86 ;
      RECT 147.95 388.06 150.33 388.56 ;
      RECT 147.95 389.46 148.55 390.7 ;
      RECT 147.95 389.76 150.33 390.26 ;
      RECT 109.46 389.46 148.55 389.76 ;
      RECT 109.46 391.96 148.55 392.26 ;
      RECT 147.95 391.02 148.55 392.26 ;
      RECT 147.95 391.46 150.33 391.96 ;
      RECT 147.95 392.86 148.55 394.1 ;
      RECT 147.95 393.16 150.33 393.66 ;
      RECT 109.46 392.86 148.55 393.16 ;
      RECT 109.46 395.36 148.55 395.66 ;
      RECT 147.95 394.42 148.55 395.66 ;
      RECT 147.95 394.86 150.33 395.36 ;
      RECT 147.95 396.26 148.55 397.5 ;
      RECT 147.95 396.56 150.33 397.06 ;
      RECT 109.46 396.26 148.55 396.56 ;
      RECT 109.46 398.76 148.55 399.06 ;
      RECT 147.95 397.82 148.55 399.06 ;
      RECT 147.95 398.26 150.33 398.76 ;
      RECT 147.95 399.66 148.55 400.9 ;
      RECT 147.95 399.96 150.33 400.46 ;
      RECT 109.46 399.66 148.55 399.96 ;
      RECT 109.46 402.16 148.55 402.46 ;
      RECT 147.95 401.22 148.55 402.46 ;
      RECT 147.95 401.66 150.33 402.16 ;
      RECT 147.95 403.06 148.55 404.3 ;
      RECT 147.95 403.36 150.33 403.86 ;
      RECT 109.46 403.06 148.55 403.36 ;
      RECT 109.46 405.56 148.55 405.86 ;
      RECT 147.95 404.62 148.55 405.86 ;
      RECT 147.95 405.06 150.33 405.56 ;
      RECT 147.95 406.46 148.55 407.7 ;
      RECT 147.95 406.76 150.33 407.26 ;
      RECT 109.46 406.46 148.55 406.76 ;
      RECT 109.46 408.96 148.55 409.26 ;
      RECT 147.95 408.02 148.55 409.26 ;
      RECT 147.95 408.46 150.33 408.96 ;
      RECT 147.95 409.86 148.55 411.1 ;
      RECT 147.95 410.16 150.33 410.66 ;
      RECT 109.46 409.86 148.55 410.16 ;
      RECT 109.46 412.36 148.55 412.66 ;
      RECT 147.95 411.42 148.55 412.66 ;
      RECT 147.95 411.86 150.33 412.36 ;
      RECT 147.95 413.26 148.55 414.5 ;
      RECT 147.95 413.56 150.33 414.06 ;
      RECT 109.46 413.26 148.55 413.56 ;
      RECT 109.46 415.76 148.55 416.06 ;
      RECT 147.95 414.82 148.55 416.06 ;
      RECT 147.95 415.26 150.33 415.76 ;
      RECT 147.95 416.66 148.55 417.9 ;
      RECT 147.95 416.96 150.33 417.46 ;
      RECT 109.46 416.66 148.55 416.96 ;
      RECT 109.46 419.16 148.55 419.46 ;
      RECT 147.95 418.22 148.55 419.46 ;
      RECT 147.95 418.66 150.33 419.16 ;
      RECT 147.95 420.06 148.55 421.3 ;
      RECT 147.95 420.36 150.33 420.86 ;
      RECT 109.46 420.06 148.55 420.36 ;
      RECT 109.46 422.56 148.55 422.86 ;
      RECT 147.95 421.62 148.55 422.86 ;
      RECT 147.95 422.06 150.33 422.56 ;
      RECT 147.95 423.46 148.55 424.7 ;
      RECT 147.95 423.76 150.33 424.26 ;
      RECT 109.46 423.46 148.55 423.76 ;
      RECT 109.46 425.96 148.55 426.26 ;
      RECT 147.95 425.02 148.55 426.26 ;
      RECT 147.95 425.46 150.33 425.96 ;
      RECT 147.95 426.86 148.55 428.1 ;
      RECT 147.95 427.16 150.33 427.66 ;
      RECT 109.46 426.86 148.55 427.16 ;
      RECT 109.46 429.36 148.55 429.66 ;
      RECT 147.95 428.42 148.55 429.66 ;
      RECT 147.95 428.86 150.33 429.36 ;
      RECT 147.95 430.26 148.55 431.5 ;
      RECT 147.95 430.56 150.33 431.06 ;
      RECT 109.46 430.26 148.55 430.56 ;
      RECT 109.46 432.76 148.55 433.06 ;
      RECT 147.95 431.82 148.55 433.06 ;
      RECT 147.95 432.26 150.33 432.76 ;
      RECT 147.95 433.66 148.55 434.9 ;
      RECT 147.95 433.96 150.33 434.46 ;
      RECT 109.46 433.66 148.55 433.96 ;
      RECT 109.46 436.16 148.55 436.46 ;
      RECT 147.95 435.22 148.55 436.46 ;
      RECT 147.95 435.66 150.33 436.16 ;
      RECT 147.95 437.06 148.55 438.3 ;
      RECT 147.95 437.36 150.33 437.86 ;
      RECT 109.46 437.06 148.55 437.36 ;
      RECT 109.46 439.56 148.55 439.86 ;
      RECT 147.95 438.62 148.55 439.86 ;
      RECT 147.95 439.06 150.33 439.56 ;
      RECT 147.95 440.46 148.55 441.7 ;
      RECT 147.95 440.76 150.33 441.26 ;
      RECT 109.46 440.46 148.55 440.76 ;
      RECT 109.46 442.96 148.55 443.26 ;
      RECT 147.95 442.02 148.55 443.26 ;
      RECT 147.95 442.46 150.33 442.96 ;
      RECT 147.95 443.86 148.55 445.1 ;
      RECT 147.95 444.16 150.33 444.66 ;
      RECT 109.46 443.86 148.55 444.16 ;
      RECT 109.46 446.36 148.55 446.66 ;
      RECT 147.95 445.42 148.55 446.66 ;
      RECT 147.95 445.86 150.33 446.36 ;
      RECT 147.95 447.26 148.55 448.5 ;
      RECT 147.95 447.56 150.33 448.06 ;
      RECT 109.46 447.26 148.55 447.56 ;
      RECT 109.46 449.76 148.55 450.06 ;
      RECT 147.95 448.82 148.55 450.06 ;
      RECT 147.95 449.26 150.33 449.76 ;
      RECT 147.95 450.66 148.55 451.9 ;
      RECT 147.95 450.96 150.33 451.46 ;
      RECT 109.46 450.66 148.55 450.96 ;
      RECT 109.46 453.16 148.55 453.46 ;
      RECT 147.95 452.22 148.55 453.46 ;
      RECT 147.95 452.66 150.33 453.16 ;
      RECT 147.95 454.06 148.55 455.3 ;
      RECT 147.95 454.36 150.33 454.86 ;
      RECT 109.46 454.06 148.55 454.36 ;
      RECT 109.46 456.56 148.55 456.86 ;
      RECT 147.95 455.62 148.55 456.86 ;
      RECT 147.95 456.06 150.33 456.56 ;
      RECT 147.95 457.46 148.55 458.7 ;
      RECT 147.95 457.76 150.33 458.26 ;
      RECT 109.46 457.46 148.55 457.76 ;
      RECT 109.46 459.96 148.55 460.26 ;
      RECT 147.95 459.02 148.55 460.26 ;
      RECT 147.95 459.46 150.33 459.96 ;
      RECT 147.95 460.86 148.55 462.1 ;
      RECT 147.95 461.16 150.33 461.66 ;
      RECT 109.46 460.86 148.55 461.16 ;
      RECT 109.46 463.36 148.55 463.66 ;
      RECT 147.95 462.42 148.55 463.66 ;
      RECT 147.95 462.86 150.33 463.36 ;
      RECT 147.95 464.26 148.55 465.5 ;
      RECT 147.95 464.56 150.33 465.06 ;
      RECT 109.46 464.26 148.55 464.56 ;
      RECT 109.46 466.76 148.55 467.06 ;
      RECT 147.95 465.82 148.55 467.06 ;
      RECT 147.95 466.26 150.33 466.76 ;
      RECT 147.95 467.66 148.55 468.9 ;
      RECT 147.95 467.96 150.33 468.46 ;
      RECT 109.46 467.66 148.55 467.96 ;
      RECT 109.46 470.16 148.55 470.46 ;
      RECT 147.95 469.22 148.55 470.46 ;
      RECT 147.95 469.66 150.33 470.16 ;
      RECT 147.95 471.06 148.55 472.3 ;
      RECT 147.95 471.36 150.33 471.86 ;
      RECT 109.46 471.06 148.55 471.36 ;
      RECT 109.46 473.56 148.55 473.86 ;
      RECT 147.95 472.62 148.55 473.86 ;
      RECT 147.95 473.06 150.33 473.56 ;
      RECT 147.95 474.46 148.55 475.7 ;
      RECT 147.95 474.76 150.33 475.26 ;
      RECT 109.46 474.46 148.55 474.76 ;
      RECT 109.46 476.96 148.55 477.26 ;
      RECT 147.95 476.02 148.55 477.26 ;
      RECT 147.95 476.46 150.33 476.96 ;
      RECT 147.95 477.86 148.55 479.1 ;
      RECT 147.95 478.16 150.33 478.66 ;
      RECT 109.46 477.86 148.55 478.16 ;
      RECT 109.46 480.36 148.55 480.66 ;
      RECT 147.95 479.42 148.55 480.66 ;
      RECT 147.95 479.86 150.33 480.36 ;
      RECT 147.95 481.26 148.55 482.5 ;
      RECT 147.95 481.56 150.33 482.06 ;
      RECT 109.46 481.26 148.55 481.56 ;
      RECT 109.46 483.76 148.55 484.06 ;
      RECT 147.95 482.82 148.55 484.06 ;
      RECT 147.95 483.26 150.33 483.76 ;
      RECT 147.95 484.66 148.55 485.9 ;
      RECT 147.95 484.96 150.33 485.46 ;
      RECT 109.46 484.66 148.55 484.96 ;
      RECT 109.46 487.16 148.55 487.46 ;
      RECT 147.95 486.22 148.55 487.46 ;
      RECT 147.95 486.66 150.33 487.16 ;
      RECT 147.95 488.06 148.55 489.3 ;
      RECT 147.95 488.36 150.33 488.86 ;
      RECT 109.46 488.06 148.55 488.36 ;
      RECT 109.46 490.56 148.55 490.86 ;
      RECT 147.95 489.62 148.55 490.86 ;
      RECT 147.95 490.06 150.33 490.56 ;
      RECT 147.95 491.46 148.55 492.7 ;
      RECT 147.95 491.76 150.33 492.26 ;
      RECT 109.46 491.46 148.55 491.76 ;
      RECT 109.46 493.96 148.55 494.26 ;
      RECT 147.95 493.02 148.55 494.26 ;
      RECT 147.95 493.46 150.33 493.96 ;
      RECT 147.95 494.86 148.55 496.1 ;
      RECT 147.95 495.16 150.33 495.66 ;
      RECT 109.46 494.86 148.55 495.16 ;
      RECT 109.46 497.36 148.55 497.66 ;
      RECT 147.95 496.42 148.55 497.66 ;
      RECT 147.95 496.86 150.33 497.36 ;
      RECT 147.95 498.26 148.55 499.5 ;
      RECT 147.95 498.56 150.33 499.06 ;
      RECT 109.46 498.26 148.55 498.56 ;
      RECT 109.46 500.76 148.55 501.06 ;
      RECT 147.95 499.82 148.55 501.06 ;
      RECT 147.95 500.26 150.33 500.76 ;
      RECT 147.95 501.66 148.55 502.9 ;
      RECT 147.95 501.96 150.33 502.46 ;
      RECT 109.46 501.66 148.55 501.96 ;
      RECT 109.46 504.16 148.55 504.46 ;
      RECT 147.95 503.22 148.55 504.46 ;
      RECT 147.95 503.66 150.33 504.16 ;
      RECT 150.13 505.14 150.33 506.9 ;
      RECT 109.46 505.14 150.33 505.34 ;
      RECT 135.4 507.58 149.01 508.1 ;
      RECT 135.4 507.58 150.01 507.78 ;
      RECT 149.01 509.8 149.79 510 ;
      RECT 149.01 508.3 149.21 510 ;
      RECT 132.41 508.3 149.21 508.5 ;
      RECT 132.41 507.22 132.61 508.5 ;
      RECT 114.94 507.22 132.61 507.42 ;
      RECT 145.66 16.67 149.47 16.87 ;
      RECT 145.66 15.95 145.86 16.87 ;
      RECT 145.34 15.95 145.86 16.15 ;
      RECT 109.39 68.43 149.33 68.63 ;
      RECT 109.39 68.13 109.99 68.63 ;
      RECT 142.11 23.26 145.85 23.46 ;
      RECT 142.11 22.99 142.31 23.46 ;
      RECT 144.01 16.14 144.67 16.34 ;
      RECT 144.01 15.74 144.21 16.34 ;
      RECT 134.98 505.94 135.89 506.14 ;
      RECT 135.69 505.82 144.62 506.02 ;
      RECT 134.98 70.9 143.22 71.1 ;
      RECT 143.02 70.66 143.22 71.1 ;
      RECT 143.02 70.66 144.2 70.86 ;
      RECT 143.02 71.66 144.2 71.86 ;
      RECT 143.02 71.42 143.22 71.86 ;
      RECT 134.98 71.42 143.22 71.62 ;
      RECT 134.98 74.3 143.22 74.5 ;
      RECT 143.02 74.06 143.22 74.5 ;
      RECT 143.02 74.06 144.2 74.26 ;
      RECT 143.02 75.06 144.2 75.26 ;
      RECT 143.02 74.82 143.22 75.26 ;
      RECT 134.98 74.82 143.22 75.02 ;
      RECT 134.98 77.7 143.22 77.9 ;
      RECT 143.02 77.46 143.22 77.9 ;
      RECT 143.02 77.46 144.2 77.66 ;
      RECT 143.02 78.46 144.2 78.66 ;
      RECT 143.02 78.22 143.22 78.66 ;
      RECT 134.98 78.22 143.22 78.42 ;
      RECT 134.98 81.1 143.22 81.3 ;
      RECT 143.02 80.86 143.22 81.3 ;
      RECT 143.02 80.86 144.2 81.06 ;
      RECT 143.02 81.86 144.2 82.06 ;
      RECT 143.02 81.62 143.22 82.06 ;
      RECT 134.98 81.62 143.22 81.82 ;
      RECT 134.98 84.5 143.22 84.7 ;
      RECT 143.02 84.26 143.22 84.7 ;
      RECT 143.02 84.26 144.2 84.46 ;
      RECT 143.02 85.26 144.2 85.46 ;
      RECT 143.02 85.02 143.22 85.46 ;
      RECT 134.98 85.02 143.22 85.22 ;
      RECT 134.98 87.9 143.22 88.1 ;
      RECT 143.02 87.66 143.22 88.1 ;
      RECT 143.02 87.66 144.2 87.86 ;
      RECT 143.02 88.66 144.2 88.86 ;
      RECT 143.02 88.42 143.22 88.86 ;
      RECT 134.98 88.42 143.22 88.62 ;
      RECT 134.98 91.3 143.22 91.5 ;
      RECT 143.02 91.06 143.22 91.5 ;
      RECT 143.02 91.06 144.2 91.26 ;
      RECT 143.02 92.06 144.2 92.26 ;
      RECT 143.02 91.82 143.22 92.26 ;
      RECT 134.98 91.82 143.22 92.02 ;
      RECT 134.98 94.7 143.22 94.9 ;
      RECT 143.02 94.46 143.22 94.9 ;
      RECT 143.02 94.46 144.2 94.66 ;
      RECT 143.02 95.46 144.2 95.66 ;
      RECT 143.02 95.22 143.22 95.66 ;
      RECT 134.98 95.22 143.22 95.42 ;
      RECT 134.98 98.1 143.22 98.3 ;
      RECT 143.02 97.86 143.22 98.3 ;
      RECT 143.02 97.86 144.2 98.06 ;
      RECT 143.02 98.86 144.2 99.06 ;
      RECT 143.02 98.62 143.22 99.06 ;
      RECT 134.98 98.62 143.22 98.82 ;
      RECT 134.98 101.5 143.22 101.7 ;
      RECT 143.02 101.26 143.22 101.7 ;
      RECT 143.02 101.26 144.2 101.46 ;
      RECT 143.02 102.26 144.2 102.46 ;
      RECT 143.02 102.02 143.22 102.46 ;
      RECT 134.98 102.02 143.22 102.22 ;
      RECT 134.98 104.9 143.22 105.1 ;
      RECT 143.02 104.66 143.22 105.1 ;
      RECT 143.02 104.66 144.2 104.86 ;
      RECT 143.02 105.66 144.2 105.86 ;
      RECT 143.02 105.42 143.22 105.86 ;
      RECT 134.98 105.42 143.22 105.62 ;
      RECT 134.98 108.3 143.22 108.5 ;
      RECT 143.02 108.06 143.22 108.5 ;
      RECT 143.02 108.06 144.2 108.26 ;
      RECT 143.02 109.06 144.2 109.26 ;
      RECT 143.02 108.82 143.22 109.26 ;
      RECT 134.98 108.82 143.22 109.02 ;
      RECT 134.98 111.7 143.22 111.9 ;
      RECT 143.02 111.46 143.22 111.9 ;
      RECT 143.02 111.46 144.2 111.66 ;
      RECT 143.02 112.46 144.2 112.66 ;
      RECT 143.02 112.22 143.22 112.66 ;
      RECT 134.98 112.22 143.22 112.42 ;
      RECT 134.98 115.1 143.22 115.3 ;
      RECT 143.02 114.86 143.22 115.3 ;
      RECT 143.02 114.86 144.2 115.06 ;
      RECT 143.02 115.86 144.2 116.06 ;
      RECT 143.02 115.62 143.22 116.06 ;
      RECT 134.98 115.62 143.22 115.82 ;
      RECT 134.98 118.5 143.22 118.7 ;
      RECT 143.02 118.26 143.22 118.7 ;
      RECT 143.02 118.26 144.2 118.46 ;
      RECT 143.02 119.26 144.2 119.46 ;
      RECT 143.02 119.02 143.22 119.46 ;
      RECT 134.98 119.02 143.22 119.22 ;
      RECT 134.98 121.9 143.22 122.1 ;
      RECT 143.02 121.66 143.22 122.1 ;
      RECT 143.02 121.66 144.2 121.86 ;
      RECT 143.02 122.66 144.2 122.86 ;
      RECT 143.02 122.42 143.22 122.86 ;
      RECT 134.98 122.42 143.22 122.62 ;
      RECT 134.98 125.3 143.22 125.5 ;
      RECT 143.02 125.06 143.22 125.5 ;
      RECT 143.02 125.06 144.2 125.26 ;
      RECT 143.02 126.06 144.2 126.26 ;
      RECT 143.02 125.82 143.22 126.26 ;
      RECT 134.98 125.82 143.22 126.02 ;
      RECT 134.98 128.7 143.22 128.9 ;
      RECT 143.02 128.46 143.22 128.9 ;
      RECT 143.02 128.46 144.2 128.66 ;
      RECT 143.02 129.46 144.2 129.66 ;
      RECT 143.02 129.22 143.22 129.66 ;
      RECT 134.98 129.22 143.22 129.42 ;
      RECT 134.98 132.1 143.22 132.3 ;
      RECT 143.02 131.86 143.22 132.3 ;
      RECT 143.02 131.86 144.2 132.06 ;
      RECT 143.02 132.86 144.2 133.06 ;
      RECT 143.02 132.62 143.22 133.06 ;
      RECT 134.98 132.62 143.22 132.82 ;
      RECT 134.98 135.5 143.22 135.7 ;
      RECT 143.02 135.26 143.22 135.7 ;
      RECT 143.02 135.26 144.2 135.46 ;
      RECT 143.02 136.26 144.2 136.46 ;
      RECT 143.02 136.02 143.22 136.46 ;
      RECT 134.98 136.02 143.22 136.22 ;
      RECT 134.98 138.9 143.22 139.1 ;
      RECT 143.02 138.66 143.22 139.1 ;
      RECT 143.02 138.66 144.2 138.86 ;
      RECT 143.02 139.66 144.2 139.86 ;
      RECT 143.02 139.42 143.22 139.86 ;
      RECT 134.98 139.42 143.22 139.62 ;
      RECT 134.98 142.3 143.22 142.5 ;
      RECT 143.02 142.06 143.22 142.5 ;
      RECT 143.02 142.06 144.2 142.26 ;
      RECT 143.02 143.06 144.2 143.26 ;
      RECT 143.02 142.82 143.22 143.26 ;
      RECT 134.98 142.82 143.22 143.02 ;
      RECT 134.98 145.7 143.22 145.9 ;
      RECT 143.02 145.46 143.22 145.9 ;
      RECT 143.02 145.46 144.2 145.66 ;
      RECT 143.02 146.46 144.2 146.66 ;
      RECT 143.02 146.22 143.22 146.66 ;
      RECT 134.98 146.22 143.22 146.42 ;
      RECT 134.98 149.1 143.22 149.3 ;
      RECT 143.02 148.86 143.22 149.3 ;
      RECT 143.02 148.86 144.2 149.06 ;
      RECT 143.02 149.86 144.2 150.06 ;
      RECT 143.02 149.62 143.22 150.06 ;
      RECT 134.98 149.62 143.22 149.82 ;
      RECT 134.98 152.5 143.22 152.7 ;
      RECT 143.02 152.26 143.22 152.7 ;
      RECT 143.02 152.26 144.2 152.46 ;
      RECT 143.02 153.26 144.2 153.46 ;
      RECT 143.02 153.02 143.22 153.46 ;
      RECT 134.98 153.02 143.22 153.22 ;
      RECT 134.98 155.9 143.22 156.1 ;
      RECT 143.02 155.66 143.22 156.1 ;
      RECT 143.02 155.66 144.2 155.86 ;
      RECT 143.02 156.66 144.2 156.86 ;
      RECT 143.02 156.42 143.22 156.86 ;
      RECT 134.98 156.42 143.22 156.62 ;
      RECT 134.98 159.3 143.22 159.5 ;
      RECT 143.02 159.06 143.22 159.5 ;
      RECT 143.02 159.06 144.2 159.26 ;
      RECT 143.02 160.06 144.2 160.26 ;
      RECT 143.02 159.82 143.22 160.26 ;
      RECT 134.98 159.82 143.22 160.02 ;
      RECT 134.98 162.7 143.22 162.9 ;
      RECT 143.02 162.46 143.22 162.9 ;
      RECT 143.02 162.46 144.2 162.66 ;
      RECT 143.02 163.46 144.2 163.66 ;
      RECT 143.02 163.22 143.22 163.66 ;
      RECT 134.98 163.22 143.22 163.42 ;
      RECT 134.98 166.1 143.22 166.3 ;
      RECT 143.02 165.86 143.22 166.3 ;
      RECT 143.02 165.86 144.2 166.06 ;
      RECT 143.02 166.86 144.2 167.06 ;
      RECT 143.02 166.62 143.22 167.06 ;
      RECT 134.98 166.62 143.22 166.82 ;
      RECT 134.98 169.5 143.22 169.7 ;
      RECT 143.02 169.26 143.22 169.7 ;
      RECT 143.02 169.26 144.2 169.46 ;
      RECT 143.02 170.26 144.2 170.46 ;
      RECT 143.02 170.02 143.22 170.46 ;
      RECT 134.98 170.02 143.22 170.22 ;
      RECT 134.98 172.9 143.22 173.1 ;
      RECT 143.02 172.66 143.22 173.1 ;
      RECT 143.02 172.66 144.2 172.86 ;
      RECT 143.02 173.66 144.2 173.86 ;
      RECT 143.02 173.42 143.22 173.86 ;
      RECT 134.98 173.42 143.22 173.62 ;
      RECT 134.98 176.3 143.22 176.5 ;
      RECT 143.02 176.06 143.22 176.5 ;
      RECT 143.02 176.06 144.2 176.26 ;
      RECT 143.02 177.06 144.2 177.26 ;
      RECT 143.02 176.82 143.22 177.26 ;
      RECT 134.98 176.82 143.22 177.02 ;
      RECT 134.98 179.7 143.22 179.9 ;
      RECT 143.02 179.46 143.22 179.9 ;
      RECT 143.02 179.46 144.2 179.66 ;
      RECT 143.02 180.46 144.2 180.66 ;
      RECT 143.02 180.22 143.22 180.66 ;
      RECT 134.98 180.22 143.22 180.42 ;
      RECT 134.98 183.1 143.22 183.3 ;
      RECT 143.02 182.86 143.22 183.3 ;
      RECT 143.02 182.86 144.2 183.06 ;
      RECT 143.02 183.86 144.2 184.06 ;
      RECT 143.02 183.62 143.22 184.06 ;
      RECT 134.98 183.62 143.22 183.82 ;
      RECT 134.98 186.5 143.22 186.7 ;
      RECT 143.02 186.26 143.22 186.7 ;
      RECT 143.02 186.26 144.2 186.46 ;
      RECT 143.02 187.26 144.2 187.46 ;
      RECT 143.02 187.02 143.22 187.46 ;
      RECT 134.98 187.02 143.22 187.22 ;
      RECT 134.98 189.9 143.22 190.1 ;
      RECT 143.02 189.66 143.22 190.1 ;
      RECT 143.02 189.66 144.2 189.86 ;
      RECT 143.02 190.66 144.2 190.86 ;
      RECT 143.02 190.42 143.22 190.86 ;
      RECT 134.98 190.42 143.22 190.62 ;
      RECT 134.98 193.3 143.22 193.5 ;
      RECT 143.02 193.06 143.22 193.5 ;
      RECT 143.02 193.06 144.2 193.26 ;
      RECT 143.02 194.06 144.2 194.26 ;
      RECT 143.02 193.82 143.22 194.26 ;
      RECT 134.98 193.82 143.22 194.02 ;
      RECT 134.98 196.7 143.22 196.9 ;
      RECT 143.02 196.46 143.22 196.9 ;
      RECT 143.02 196.46 144.2 196.66 ;
      RECT 143.02 197.46 144.2 197.66 ;
      RECT 143.02 197.22 143.22 197.66 ;
      RECT 134.98 197.22 143.22 197.42 ;
      RECT 134.98 200.1 143.22 200.3 ;
      RECT 143.02 199.86 143.22 200.3 ;
      RECT 143.02 199.86 144.2 200.06 ;
      RECT 143.02 200.86 144.2 201.06 ;
      RECT 143.02 200.62 143.22 201.06 ;
      RECT 134.98 200.62 143.22 200.82 ;
      RECT 134.98 203.5 143.22 203.7 ;
      RECT 143.02 203.26 143.22 203.7 ;
      RECT 143.02 203.26 144.2 203.46 ;
      RECT 143.02 204.26 144.2 204.46 ;
      RECT 143.02 204.02 143.22 204.46 ;
      RECT 134.98 204.02 143.22 204.22 ;
      RECT 134.98 206.9 143.22 207.1 ;
      RECT 143.02 206.66 143.22 207.1 ;
      RECT 143.02 206.66 144.2 206.86 ;
      RECT 143.02 207.66 144.2 207.86 ;
      RECT 143.02 207.42 143.22 207.86 ;
      RECT 134.98 207.42 143.22 207.62 ;
      RECT 134.98 210.3 143.22 210.5 ;
      RECT 143.02 210.06 143.22 210.5 ;
      RECT 143.02 210.06 144.2 210.26 ;
      RECT 143.02 211.06 144.2 211.26 ;
      RECT 143.02 210.82 143.22 211.26 ;
      RECT 134.98 210.82 143.22 211.02 ;
      RECT 134.98 213.7 143.22 213.9 ;
      RECT 143.02 213.46 143.22 213.9 ;
      RECT 143.02 213.46 144.2 213.66 ;
      RECT 143.02 214.46 144.2 214.66 ;
      RECT 143.02 214.22 143.22 214.66 ;
      RECT 134.98 214.22 143.22 214.42 ;
      RECT 134.98 217.1 143.22 217.3 ;
      RECT 143.02 216.86 143.22 217.3 ;
      RECT 143.02 216.86 144.2 217.06 ;
      RECT 143.02 217.86 144.2 218.06 ;
      RECT 143.02 217.62 143.22 218.06 ;
      RECT 134.98 217.62 143.22 217.82 ;
      RECT 134.98 220.5 143.22 220.7 ;
      RECT 143.02 220.26 143.22 220.7 ;
      RECT 143.02 220.26 144.2 220.46 ;
      RECT 143.02 221.26 144.2 221.46 ;
      RECT 143.02 221.02 143.22 221.46 ;
      RECT 134.98 221.02 143.22 221.22 ;
      RECT 134.98 223.9 143.22 224.1 ;
      RECT 143.02 223.66 143.22 224.1 ;
      RECT 143.02 223.66 144.2 223.86 ;
      RECT 143.02 224.66 144.2 224.86 ;
      RECT 143.02 224.42 143.22 224.86 ;
      RECT 134.98 224.42 143.22 224.62 ;
      RECT 134.98 227.3 143.22 227.5 ;
      RECT 143.02 227.06 143.22 227.5 ;
      RECT 143.02 227.06 144.2 227.26 ;
      RECT 143.02 228.06 144.2 228.26 ;
      RECT 143.02 227.82 143.22 228.26 ;
      RECT 134.98 227.82 143.22 228.02 ;
      RECT 134.98 230.7 143.22 230.9 ;
      RECT 143.02 230.46 143.22 230.9 ;
      RECT 143.02 230.46 144.2 230.66 ;
      RECT 143.02 231.46 144.2 231.66 ;
      RECT 143.02 231.22 143.22 231.66 ;
      RECT 134.98 231.22 143.22 231.42 ;
      RECT 134.98 234.1 143.22 234.3 ;
      RECT 143.02 233.86 143.22 234.3 ;
      RECT 143.02 233.86 144.2 234.06 ;
      RECT 143.02 234.86 144.2 235.06 ;
      RECT 143.02 234.62 143.22 235.06 ;
      RECT 134.98 234.62 143.22 234.82 ;
      RECT 134.98 237.5 143.22 237.7 ;
      RECT 143.02 237.26 143.22 237.7 ;
      RECT 143.02 237.26 144.2 237.46 ;
      RECT 143.02 238.26 144.2 238.46 ;
      RECT 143.02 238.02 143.22 238.46 ;
      RECT 134.98 238.02 143.22 238.22 ;
      RECT 134.98 240.9 143.22 241.1 ;
      RECT 143.02 240.66 143.22 241.1 ;
      RECT 143.02 240.66 144.2 240.86 ;
      RECT 143.02 241.66 144.2 241.86 ;
      RECT 143.02 241.42 143.22 241.86 ;
      RECT 134.98 241.42 143.22 241.62 ;
      RECT 134.98 244.3 143.22 244.5 ;
      RECT 143.02 244.06 143.22 244.5 ;
      RECT 143.02 244.06 144.2 244.26 ;
      RECT 143.02 245.06 144.2 245.26 ;
      RECT 143.02 244.82 143.22 245.26 ;
      RECT 134.98 244.82 143.22 245.02 ;
      RECT 134.98 247.7 143.22 247.9 ;
      RECT 143.02 247.46 143.22 247.9 ;
      RECT 143.02 247.46 144.2 247.66 ;
      RECT 143.02 248.46 144.2 248.66 ;
      RECT 143.02 248.22 143.22 248.66 ;
      RECT 134.98 248.22 143.22 248.42 ;
      RECT 134.98 251.1 143.22 251.3 ;
      RECT 143.02 250.86 143.22 251.3 ;
      RECT 143.02 250.86 144.2 251.06 ;
      RECT 143.02 251.86 144.2 252.06 ;
      RECT 143.02 251.62 143.22 252.06 ;
      RECT 134.98 251.62 143.22 251.82 ;
      RECT 134.98 254.5 143.22 254.7 ;
      RECT 143.02 254.26 143.22 254.7 ;
      RECT 143.02 254.26 144.2 254.46 ;
      RECT 143.02 255.26 144.2 255.46 ;
      RECT 143.02 255.02 143.22 255.46 ;
      RECT 134.98 255.02 143.22 255.22 ;
      RECT 134.98 257.9 143.22 258.1 ;
      RECT 143.02 257.66 143.22 258.1 ;
      RECT 143.02 257.66 144.2 257.86 ;
      RECT 143.02 258.66 144.2 258.86 ;
      RECT 143.02 258.42 143.22 258.86 ;
      RECT 134.98 258.42 143.22 258.62 ;
      RECT 134.98 261.3 143.22 261.5 ;
      RECT 143.02 261.06 143.22 261.5 ;
      RECT 143.02 261.06 144.2 261.26 ;
      RECT 143.02 262.06 144.2 262.26 ;
      RECT 143.02 261.82 143.22 262.26 ;
      RECT 134.98 261.82 143.22 262.02 ;
      RECT 134.98 264.7 143.22 264.9 ;
      RECT 143.02 264.46 143.22 264.9 ;
      RECT 143.02 264.46 144.2 264.66 ;
      RECT 143.02 265.46 144.2 265.66 ;
      RECT 143.02 265.22 143.22 265.66 ;
      RECT 134.98 265.22 143.22 265.42 ;
      RECT 134.98 268.1 143.22 268.3 ;
      RECT 143.02 267.86 143.22 268.3 ;
      RECT 143.02 267.86 144.2 268.06 ;
      RECT 143.02 268.86 144.2 269.06 ;
      RECT 143.02 268.62 143.22 269.06 ;
      RECT 134.98 268.62 143.22 268.82 ;
      RECT 134.98 271.5 143.22 271.7 ;
      RECT 143.02 271.26 143.22 271.7 ;
      RECT 143.02 271.26 144.2 271.46 ;
      RECT 143.02 272.26 144.2 272.46 ;
      RECT 143.02 272.02 143.22 272.46 ;
      RECT 134.98 272.02 143.22 272.22 ;
      RECT 134.98 274.9 143.22 275.1 ;
      RECT 143.02 274.66 143.22 275.1 ;
      RECT 143.02 274.66 144.2 274.86 ;
      RECT 143.02 275.66 144.2 275.86 ;
      RECT 143.02 275.42 143.22 275.86 ;
      RECT 134.98 275.42 143.22 275.62 ;
      RECT 134.98 278.3 143.22 278.5 ;
      RECT 143.02 278.06 143.22 278.5 ;
      RECT 143.02 278.06 144.2 278.26 ;
      RECT 143.02 279.06 144.2 279.26 ;
      RECT 143.02 278.82 143.22 279.26 ;
      RECT 134.98 278.82 143.22 279.02 ;
      RECT 134.98 281.7 143.22 281.9 ;
      RECT 143.02 281.46 143.22 281.9 ;
      RECT 143.02 281.46 144.2 281.66 ;
      RECT 143.02 282.46 144.2 282.66 ;
      RECT 143.02 282.22 143.22 282.66 ;
      RECT 134.98 282.22 143.22 282.42 ;
      RECT 134.98 285.1 143.22 285.3 ;
      RECT 143.02 284.86 143.22 285.3 ;
      RECT 143.02 284.86 144.2 285.06 ;
      RECT 143.02 285.86 144.2 286.06 ;
      RECT 143.02 285.62 143.22 286.06 ;
      RECT 134.98 285.62 143.22 285.82 ;
      RECT 134.98 288.5 143.22 288.7 ;
      RECT 143.02 288.26 143.22 288.7 ;
      RECT 143.02 288.26 144.2 288.46 ;
      RECT 143.02 289.26 144.2 289.46 ;
      RECT 143.02 289.02 143.22 289.46 ;
      RECT 134.98 289.02 143.22 289.22 ;
      RECT 134.98 291.9 143.22 292.1 ;
      RECT 143.02 291.66 143.22 292.1 ;
      RECT 143.02 291.66 144.2 291.86 ;
      RECT 143.02 292.66 144.2 292.86 ;
      RECT 143.02 292.42 143.22 292.86 ;
      RECT 134.98 292.42 143.22 292.62 ;
      RECT 134.98 295.3 143.22 295.5 ;
      RECT 143.02 295.06 143.22 295.5 ;
      RECT 143.02 295.06 144.2 295.26 ;
      RECT 143.02 296.06 144.2 296.26 ;
      RECT 143.02 295.82 143.22 296.26 ;
      RECT 134.98 295.82 143.22 296.02 ;
      RECT 134.98 298.7 143.22 298.9 ;
      RECT 143.02 298.46 143.22 298.9 ;
      RECT 143.02 298.46 144.2 298.66 ;
      RECT 143.02 299.46 144.2 299.66 ;
      RECT 143.02 299.22 143.22 299.66 ;
      RECT 134.98 299.22 143.22 299.42 ;
      RECT 134.98 302.1 143.22 302.3 ;
      RECT 143.02 301.86 143.22 302.3 ;
      RECT 143.02 301.86 144.2 302.06 ;
      RECT 143.02 302.86 144.2 303.06 ;
      RECT 143.02 302.62 143.22 303.06 ;
      RECT 134.98 302.62 143.22 302.82 ;
      RECT 134.98 305.5 143.22 305.7 ;
      RECT 143.02 305.26 143.22 305.7 ;
      RECT 143.02 305.26 144.2 305.46 ;
      RECT 143.02 306.26 144.2 306.46 ;
      RECT 143.02 306.02 143.22 306.46 ;
      RECT 134.98 306.02 143.22 306.22 ;
      RECT 134.98 308.9 143.22 309.1 ;
      RECT 143.02 308.66 143.22 309.1 ;
      RECT 143.02 308.66 144.2 308.86 ;
      RECT 143.02 309.66 144.2 309.86 ;
      RECT 143.02 309.42 143.22 309.86 ;
      RECT 134.98 309.42 143.22 309.62 ;
      RECT 134.98 312.3 143.22 312.5 ;
      RECT 143.02 312.06 143.22 312.5 ;
      RECT 143.02 312.06 144.2 312.26 ;
      RECT 143.02 313.06 144.2 313.26 ;
      RECT 143.02 312.82 143.22 313.26 ;
      RECT 134.98 312.82 143.22 313.02 ;
      RECT 134.98 315.7 143.22 315.9 ;
      RECT 143.02 315.46 143.22 315.9 ;
      RECT 143.02 315.46 144.2 315.66 ;
      RECT 143.02 316.46 144.2 316.66 ;
      RECT 143.02 316.22 143.22 316.66 ;
      RECT 134.98 316.22 143.22 316.42 ;
      RECT 134.98 319.1 143.22 319.3 ;
      RECT 143.02 318.86 143.22 319.3 ;
      RECT 143.02 318.86 144.2 319.06 ;
      RECT 143.02 319.86 144.2 320.06 ;
      RECT 143.02 319.62 143.22 320.06 ;
      RECT 134.98 319.62 143.22 319.82 ;
      RECT 134.98 322.5 143.22 322.7 ;
      RECT 143.02 322.26 143.22 322.7 ;
      RECT 143.02 322.26 144.2 322.46 ;
      RECT 143.02 323.26 144.2 323.46 ;
      RECT 143.02 323.02 143.22 323.46 ;
      RECT 134.98 323.02 143.22 323.22 ;
      RECT 134.98 325.9 143.22 326.1 ;
      RECT 143.02 325.66 143.22 326.1 ;
      RECT 143.02 325.66 144.2 325.86 ;
      RECT 143.02 326.66 144.2 326.86 ;
      RECT 143.02 326.42 143.22 326.86 ;
      RECT 134.98 326.42 143.22 326.62 ;
      RECT 134.98 329.3 143.22 329.5 ;
      RECT 143.02 329.06 143.22 329.5 ;
      RECT 143.02 329.06 144.2 329.26 ;
      RECT 143.02 330.06 144.2 330.26 ;
      RECT 143.02 329.82 143.22 330.26 ;
      RECT 134.98 329.82 143.22 330.02 ;
      RECT 134.98 332.7 143.22 332.9 ;
      RECT 143.02 332.46 143.22 332.9 ;
      RECT 143.02 332.46 144.2 332.66 ;
      RECT 143.02 333.46 144.2 333.66 ;
      RECT 143.02 333.22 143.22 333.66 ;
      RECT 134.98 333.22 143.22 333.42 ;
      RECT 134.98 336.1 143.22 336.3 ;
      RECT 143.02 335.86 143.22 336.3 ;
      RECT 143.02 335.86 144.2 336.06 ;
      RECT 143.02 336.86 144.2 337.06 ;
      RECT 143.02 336.62 143.22 337.06 ;
      RECT 134.98 336.62 143.22 336.82 ;
      RECT 134.98 339.5 143.22 339.7 ;
      RECT 143.02 339.26 143.22 339.7 ;
      RECT 143.02 339.26 144.2 339.46 ;
      RECT 143.02 340.26 144.2 340.46 ;
      RECT 143.02 340.02 143.22 340.46 ;
      RECT 134.98 340.02 143.22 340.22 ;
      RECT 134.98 342.9 143.22 343.1 ;
      RECT 143.02 342.66 143.22 343.1 ;
      RECT 143.02 342.66 144.2 342.86 ;
      RECT 143.02 343.66 144.2 343.86 ;
      RECT 143.02 343.42 143.22 343.86 ;
      RECT 134.98 343.42 143.22 343.62 ;
      RECT 134.98 346.3 143.22 346.5 ;
      RECT 143.02 346.06 143.22 346.5 ;
      RECT 143.02 346.06 144.2 346.26 ;
      RECT 143.02 347.06 144.2 347.26 ;
      RECT 143.02 346.82 143.22 347.26 ;
      RECT 134.98 346.82 143.22 347.02 ;
      RECT 134.98 349.7 143.22 349.9 ;
      RECT 143.02 349.46 143.22 349.9 ;
      RECT 143.02 349.46 144.2 349.66 ;
      RECT 143.02 350.46 144.2 350.66 ;
      RECT 143.02 350.22 143.22 350.66 ;
      RECT 134.98 350.22 143.22 350.42 ;
      RECT 134.98 353.1 143.22 353.3 ;
      RECT 143.02 352.86 143.22 353.3 ;
      RECT 143.02 352.86 144.2 353.06 ;
      RECT 143.02 353.86 144.2 354.06 ;
      RECT 143.02 353.62 143.22 354.06 ;
      RECT 134.98 353.62 143.22 353.82 ;
      RECT 134.98 356.5 143.22 356.7 ;
      RECT 143.02 356.26 143.22 356.7 ;
      RECT 143.02 356.26 144.2 356.46 ;
      RECT 143.02 357.26 144.2 357.46 ;
      RECT 143.02 357.02 143.22 357.46 ;
      RECT 134.98 357.02 143.22 357.22 ;
      RECT 134.98 359.9 143.22 360.1 ;
      RECT 143.02 359.66 143.22 360.1 ;
      RECT 143.02 359.66 144.2 359.86 ;
      RECT 143.02 360.66 144.2 360.86 ;
      RECT 143.02 360.42 143.22 360.86 ;
      RECT 134.98 360.42 143.22 360.62 ;
      RECT 134.98 363.3 143.22 363.5 ;
      RECT 143.02 363.06 143.22 363.5 ;
      RECT 143.02 363.06 144.2 363.26 ;
      RECT 143.02 364.06 144.2 364.26 ;
      RECT 143.02 363.82 143.22 364.26 ;
      RECT 134.98 363.82 143.22 364.02 ;
      RECT 134.98 366.7 143.22 366.9 ;
      RECT 143.02 366.46 143.22 366.9 ;
      RECT 143.02 366.46 144.2 366.66 ;
      RECT 143.02 367.46 144.2 367.66 ;
      RECT 143.02 367.22 143.22 367.66 ;
      RECT 134.98 367.22 143.22 367.42 ;
      RECT 134.98 370.1 143.22 370.3 ;
      RECT 143.02 369.86 143.22 370.3 ;
      RECT 143.02 369.86 144.2 370.06 ;
      RECT 143.02 370.86 144.2 371.06 ;
      RECT 143.02 370.62 143.22 371.06 ;
      RECT 134.98 370.62 143.22 370.82 ;
      RECT 134.98 373.5 143.22 373.7 ;
      RECT 143.02 373.26 143.22 373.7 ;
      RECT 143.02 373.26 144.2 373.46 ;
      RECT 143.02 374.26 144.2 374.46 ;
      RECT 143.02 374.02 143.22 374.46 ;
      RECT 134.98 374.02 143.22 374.22 ;
      RECT 134.98 376.9 143.22 377.1 ;
      RECT 143.02 376.66 143.22 377.1 ;
      RECT 143.02 376.66 144.2 376.86 ;
      RECT 143.02 377.66 144.2 377.86 ;
      RECT 143.02 377.42 143.22 377.86 ;
      RECT 134.98 377.42 143.22 377.62 ;
      RECT 134.98 380.3 143.22 380.5 ;
      RECT 143.02 380.06 143.22 380.5 ;
      RECT 143.02 380.06 144.2 380.26 ;
      RECT 143.02 381.06 144.2 381.26 ;
      RECT 143.02 380.82 143.22 381.26 ;
      RECT 134.98 380.82 143.22 381.02 ;
      RECT 134.98 383.7 143.22 383.9 ;
      RECT 143.02 383.46 143.22 383.9 ;
      RECT 143.02 383.46 144.2 383.66 ;
      RECT 143.02 384.46 144.2 384.66 ;
      RECT 143.02 384.22 143.22 384.66 ;
      RECT 134.98 384.22 143.22 384.42 ;
      RECT 134.98 387.1 143.22 387.3 ;
      RECT 143.02 386.86 143.22 387.3 ;
      RECT 143.02 386.86 144.2 387.06 ;
      RECT 143.02 387.86 144.2 388.06 ;
      RECT 143.02 387.62 143.22 388.06 ;
      RECT 134.98 387.62 143.22 387.82 ;
      RECT 134.98 390.5 143.22 390.7 ;
      RECT 143.02 390.26 143.22 390.7 ;
      RECT 143.02 390.26 144.2 390.46 ;
      RECT 143.02 391.26 144.2 391.46 ;
      RECT 143.02 391.02 143.22 391.46 ;
      RECT 134.98 391.02 143.22 391.22 ;
      RECT 134.98 393.9 143.22 394.1 ;
      RECT 143.02 393.66 143.22 394.1 ;
      RECT 143.02 393.66 144.2 393.86 ;
      RECT 143.02 394.66 144.2 394.86 ;
      RECT 143.02 394.42 143.22 394.86 ;
      RECT 134.98 394.42 143.22 394.62 ;
      RECT 134.98 397.3 143.22 397.5 ;
      RECT 143.02 397.06 143.22 397.5 ;
      RECT 143.02 397.06 144.2 397.26 ;
      RECT 143.02 398.06 144.2 398.26 ;
      RECT 143.02 397.82 143.22 398.26 ;
      RECT 134.98 397.82 143.22 398.02 ;
      RECT 134.98 400.7 143.22 400.9 ;
      RECT 143.02 400.46 143.22 400.9 ;
      RECT 143.02 400.46 144.2 400.66 ;
      RECT 143.02 401.46 144.2 401.66 ;
      RECT 143.02 401.22 143.22 401.66 ;
      RECT 134.98 401.22 143.22 401.42 ;
      RECT 134.98 404.1 143.22 404.3 ;
      RECT 143.02 403.86 143.22 404.3 ;
      RECT 143.02 403.86 144.2 404.06 ;
      RECT 143.02 404.86 144.2 405.06 ;
      RECT 143.02 404.62 143.22 405.06 ;
      RECT 134.98 404.62 143.22 404.82 ;
      RECT 134.98 407.5 143.22 407.7 ;
      RECT 143.02 407.26 143.22 407.7 ;
      RECT 143.02 407.26 144.2 407.46 ;
      RECT 143.02 408.26 144.2 408.46 ;
      RECT 143.02 408.02 143.22 408.46 ;
      RECT 134.98 408.02 143.22 408.22 ;
      RECT 134.98 410.9 143.22 411.1 ;
      RECT 143.02 410.66 143.22 411.1 ;
      RECT 143.02 410.66 144.2 410.86 ;
      RECT 143.02 411.66 144.2 411.86 ;
      RECT 143.02 411.42 143.22 411.86 ;
      RECT 134.98 411.42 143.22 411.62 ;
      RECT 134.98 414.3 143.22 414.5 ;
      RECT 143.02 414.06 143.22 414.5 ;
      RECT 143.02 414.06 144.2 414.26 ;
      RECT 143.02 415.06 144.2 415.26 ;
      RECT 143.02 414.82 143.22 415.26 ;
      RECT 134.98 414.82 143.22 415.02 ;
      RECT 134.98 417.7 143.22 417.9 ;
      RECT 143.02 417.46 143.22 417.9 ;
      RECT 143.02 417.46 144.2 417.66 ;
      RECT 143.02 418.46 144.2 418.66 ;
      RECT 143.02 418.22 143.22 418.66 ;
      RECT 134.98 418.22 143.22 418.42 ;
      RECT 134.98 421.1 143.22 421.3 ;
      RECT 143.02 420.86 143.22 421.3 ;
      RECT 143.02 420.86 144.2 421.06 ;
      RECT 143.02 421.86 144.2 422.06 ;
      RECT 143.02 421.62 143.22 422.06 ;
      RECT 134.98 421.62 143.22 421.82 ;
      RECT 134.98 424.5 143.22 424.7 ;
      RECT 143.02 424.26 143.22 424.7 ;
      RECT 143.02 424.26 144.2 424.46 ;
      RECT 143.02 425.26 144.2 425.46 ;
      RECT 143.02 425.02 143.22 425.46 ;
      RECT 134.98 425.02 143.22 425.22 ;
      RECT 134.98 427.9 143.22 428.1 ;
      RECT 143.02 427.66 143.22 428.1 ;
      RECT 143.02 427.66 144.2 427.86 ;
      RECT 143.02 428.66 144.2 428.86 ;
      RECT 143.02 428.42 143.22 428.86 ;
      RECT 134.98 428.42 143.22 428.62 ;
      RECT 134.98 431.3 143.22 431.5 ;
      RECT 143.02 431.06 143.22 431.5 ;
      RECT 143.02 431.06 144.2 431.26 ;
      RECT 143.02 432.06 144.2 432.26 ;
      RECT 143.02 431.82 143.22 432.26 ;
      RECT 134.98 431.82 143.22 432.02 ;
      RECT 134.98 434.7 143.22 434.9 ;
      RECT 143.02 434.46 143.22 434.9 ;
      RECT 143.02 434.46 144.2 434.66 ;
      RECT 143.02 435.46 144.2 435.66 ;
      RECT 143.02 435.22 143.22 435.66 ;
      RECT 134.98 435.22 143.22 435.42 ;
      RECT 134.98 438.1 143.22 438.3 ;
      RECT 143.02 437.86 143.22 438.3 ;
      RECT 143.02 437.86 144.2 438.06 ;
      RECT 143.02 438.86 144.2 439.06 ;
      RECT 143.02 438.62 143.22 439.06 ;
      RECT 134.98 438.62 143.22 438.82 ;
      RECT 134.98 441.5 143.22 441.7 ;
      RECT 143.02 441.26 143.22 441.7 ;
      RECT 143.02 441.26 144.2 441.46 ;
      RECT 143.02 442.26 144.2 442.46 ;
      RECT 143.02 442.02 143.22 442.46 ;
      RECT 134.98 442.02 143.22 442.22 ;
      RECT 134.98 444.9 143.22 445.1 ;
      RECT 143.02 444.66 143.22 445.1 ;
      RECT 143.02 444.66 144.2 444.86 ;
      RECT 143.02 445.66 144.2 445.86 ;
      RECT 143.02 445.42 143.22 445.86 ;
      RECT 134.98 445.42 143.22 445.62 ;
      RECT 134.98 448.3 143.22 448.5 ;
      RECT 143.02 448.06 143.22 448.5 ;
      RECT 143.02 448.06 144.2 448.26 ;
      RECT 143.02 449.06 144.2 449.26 ;
      RECT 143.02 448.82 143.22 449.26 ;
      RECT 134.98 448.82 143.22 449.02 ;
      RECT 134.98 451.7 143.22 451.9 ;
      RECT 143.02 451.46 143.22 451.9 ;
      RECT 143.02 451.46 144.2 451.66 ;
      RECT 143.02 452.46 144.2 452.66 ;
      RECT 143.02 452.22 143.22 452.66 ;
      RECT 134.98 452.22 143.22 452.42 ;
      RECT 134.98 455.1 143.22 455.3 ;
      RECT 143.02 454.86 143.22 455.3 ;
      RECT 143.02 454.86 144.2 455.06 ;
      RECT 143.02 455.86 144.2 456.06 ;
      RECT 143.02 455.62 143.22 456.06 ;
      RECT 134.98 455.62 143.22 455.82 ;
      RECT 134.98 458.5 143.22 458.7 ;
      RECT 143.02 458.26 143.22 458.7 ;
      RECT 143.02 458.26 144.2 458.46 ;
      RECT 143.02 459.26 144.2 459.46 ;
      RECT 143.02 459.02 143.22 459.46 ;
      RECT 134.98 459.02 143.22 459.22 ;
      RECT 134.98 461.9 143.22 462.1 ;
      RECT 143.02 461.66 143.22 462.1 ;
      RECT 143.02 461.66 144.2 461.86 ;
      RECT 143.02 462.66 144.2 462.86 ;
      RECT 143.02 462.42 143.22 462.86 ;
      RECT 134.98 462.42 143.22 462.62 ;
      RECT 134.98 465.3 143.22 465.5 ;
      RECT 143.02 465.06 143.22 465.5 ;
      RECT 143.02 465.06 144.2 465.26 ;
      RECT 143.02 466.06 144.2 466.26 ;
      RECT 143.02 465.82 143.22 466.26 ;
      RECT 134.98 465.82 143.22 466.02 ;
      RECT 134.98 468.7 143.22 468.9 ;
      RECT 143.02 468.46 143.22 468.9 ;
      RECT 143.02 468.46 144.2 468.66 ;
      RECT 143.02 469.46 144.2 469.66 ;
      RECT 143.02 469.22 143.22 469.66 ;
      RECT 134.98 469.22 143.22 469.42 ;
      RECT 134.98 472.1 143.22 472.3 ;
      RECT 143.02 471.86 143.22 472.3 ;
      RECT 143.02 471.86 144.2 472.06 ;
      RECT 143.02 472.86 144.2 473.06 ;
      RECT 143.02 472.62 143.22 473.06 ;
      RECT 134.98 472.62 143.22 472.82 ;
      RECT 134.98 475.5 143.22 475.7 ;
      RECT 143.02 475.26 143.22 475.7 ;
      RECT 143.02 475.26 144.2 475.46 ;
      RECT 143.02 476.26 144.2 476.46 ;
      RECT 143.02 476.02 143.22 476.46 ;
      RECT 134.98 476.02 143.22 476.22 ;
      RECT 134.98 478.9 143.22 479.1 ;
      RECT 143.02 478.66 143.22 479.1 ;
      RECT 143.02 478.66 144.2 478.86 ;
      RECT 143.02 479.66 144.2 479.86 ;
      RECT 143.02 479.42 143.22 479.86 ;
      RECT 134.98 479.42 143.22 479.62 ;
      RECT 134.98 482.3 143.22 482.5 ;
      RECT 143.02 482.06 143.22 482.5 ;
      RECT 143.02 482.06 144.2 482.26 ;
      RECT 143.02 483.06 144.2 483.26 ;
      RECT 143.02 482.82 143.22 483.26 ;
      RECT 134.98 482.82 143.22 483.02 ;
      RECT 134.98 485.7 143.22 485.9 ;
      RECT 143.02 485.46 143.22 485.9 ;
      RECT 143.02 485.46 144.2 485.66 ;
      RECT 143.02 486.46 144.2 486.66 ;
      RECT 143.02 486.22 143.22 486.66 ;
      RECT 134.98 486.22 143.22 486.42 ;
      RECT 134.98 489.1 143.22 489.3 ;
      RECT 143.02 488.86 143.22 489.3 ;
      RECT 143.02 488.86 144.2 489.06 ;
      RECT 143.02 489.86 144.2 490.06 ;
      RECT 143.02 489.62 143.22 490.06 ;
      RECT 134.98 489.62 143.22 489.82 ;
      RECT 134.98 492.5 143.22 492.7 ;
      RECT 143.02 492.26 143.22 492.7 ;
      RECT 143.02 492.26 144.2 492.46 ;
      RECT 143.02 493.26 144.2 493.46 ;
      RECT 143.02 493.02 143.22 493.46 ;
      RECT 134.98 493.02 143.22 493.22 ;
      RECT 134.98 495.9 143.22 496.1 ;
      RECT 143.02 495.66 143.22 496.1 ;
      RECT 143.02 495.66 144.2 495.86 ;
      RECT 143.02 496.66 144.2 496.86 ;
      RECT 143.02 496.42 143.22 496.86 ;
      RECT 134.98 496.42 143.22 496.62 ;
      RECT 134.98 499.3 143.22 499.5 ;
      RECT 143.02 499.06 143.22 499.5 ;
      RECT 143.02 499.06 144.2 499.26 ;
      RECT 143.02 500.06 144.2 500.26 ;
      RECT 143.02 499.82 143.22 500.26 ;
      RECT 134.98 499.82 143.22 500.02 ;
      RECT 134.98 502.7 143.22 502.9 ;
      RECT 143.02 502.46 143.22 502.9 ;
      RECT 143.02 502.46 144.2 502.66 ;
      RECT 143.02 503.46 144.2 503.66 ;
      RECT 143.02 503.22 143.22 503.66 ;
      RECT 134.98 503.22 143.22 503.42 ;
      RECT 141.43 65.83 142.47 66.63 ;
      RECT 140.21 65.83 142.47 66.23 ;
      RECT 133.81 506.34 136.95 506.54 ;
      RECT 133.81 505.54 134.01 506.54 ;
      RECT 122.82 505.54 134.01 505.74 ;
      RECT 135.62 37.14 135.82 38.38 ;
      RECT 130.2 37.14 130.4 38.38 ;
      RECT 130.2 37.14 135.82 37.34 ;
      RECT 123.81 38.64 135.41 39.08 ;
      RECT 135.01 37.58 135.41 39.08 ;
      RECT 128.21 38.62 135.41 39.08 ;
      RECT 123.81 37.58 124.21 39.08 ;
      RECT 130.61 37.58 131.01 39.08 ;
      RECT 128.21 37.58 128.61 39.08 ;
      RECT 126.68 70.76 130.12 70.96 ;
      RECT 129.92 70.66 130.52 70.86 ;
      RECT 129.92 71.66 130.52 71.86 ;
      RECT 126.68 71.56 130.12 71.76 ;
      RECT 126.68 74.16 130.12 74.36 ;
      RECT 129.92 74.06 130.52 74.26 ;
      RECT 129.92 75.06 130.52 75.26 ;
      RECT 126.68 74.96 130.12 75.16 ;
      RECT 126.68 77.56 130.12 77.76 ;
      RECT 129.92 77.46 130.52 77.66 ;
      RECT 129.92 78.46 130.52 78.66 ;
      RECT 126.68 78.36 130.12 78.56 ;
      RECT 126.68 80.96 130.12 81.16 ;
      RECT 129.92 80.86 130.52 81.06 ;
      RECT 129.92 81.86 130.52 82.06 ;
      RECT 126.68 81.76 130.12 81.96 ;
      RECT 126.68 84.36 130.12 84.56 ;
      RECT 129.92 84.26 130.52 84.46 ;
      RECT 129.92 85.26 130.52 85.46 ;
      RECT 126.68 85.16 130.12 85.36 ;
      RECT 126.68 87.76 130.12 87.96 ;
      RECT 129.92 87.66 130.52 87.86 ;
      RECT 129.92 88.66 130.52 88.86 ;
      RECT 126.68 88.56 130.12 88.76 ;
      RECT 126.68 91.16 130.12 91.36 ;
      RECT 129.92 91.06 130.52 91.26 ;
      RECT 129.92 92.06 130.52 92.26 ;
      RECT 126.68 91.96 130.12 92.16 ;
      RECT 126.68 94.56 130.12 94.76 ;
      RECT 129.92 94.46 130.52 94.66 ;
      RECT 129.92 95.46 130.52 95.66 ;
      RECT 126.68 95.36 130.12 95.56 ;
      RECT 126.68 97.96 130.12 98.16 ;
      RECT 129.92 97.86 130.52 98.06 ;
      RECT 129.92 98.86 130.52 99.06 ;
      RECT 126.68 98.76 130.12 98.96 ;
      RECT 126.68 101.36 130.12 101.56 ;
      RECT 129.92 101.26 130.52 101.46 ;
      RECT 129.92 102.26 130.52 102.46 ;
      RECT 126.68 102.16 130.12 102.36 ;
      RECT 126.68 104.76 130.12 104.96 ;
      RECT 129.92 104.66 130.52 104.86 ;
      RECT 129.92 105.66 130.52 105.86 ;
      RECT 126.68 105.56 130.12 105.76 ;
      RECT 126.68 108.16 130.12 108.36 ;
      RECT 129.92 108.06 130.52 108.26 ;
      RECT 129.92 109.06 130.52 109.26 ;
      RECT 126.68 108.96 130.12 109.16 ;
      RECT 126.68 111.56 130.12 111.76 ;
      RECT 129.92 111.46 130.52 111.66 ;
      RECT 129.92 112.46 130.52 112.66 ;
      RECT 126.68 112.36 130.12 112.56 ;
      RECT 126.68 114.96 130.12 115.16 ;
      RECT 129.92 114.86 130.52 115.06 ;
      RECT 129.92 115.86 130.52 116.06 ;
      RECT 126.68 115.76 130.12 115.96 ;
      RECT 126.68 118.36 130.12 118.56 ;
      RECT 129.92 118.26 130.52 118.46 ;
      RECT 129.92 119.26 130.52 119.46 ;
      RECT 126.68 119.16 130.12 119.36 ;
      RECT 126.68 121.76 130.12 121.96 ;
      RECT 129.92 121.66 130.52 121.86 ;
      RECT 129.92 122.66 130.52 122.86 ;
      RECT 126.68 122.56 130.12 122.76 ;
      RECT 126.68 125.16 130.12 125.36 ;
      RECT 129.92 125.06 130.52 125.26 ;
      RECT 129.92 126.06 130.52 126.26 ;
      RECT 126.68 125.96 130.12 126.16 ;
      RECT 126.68 128.56 130.12 128.76 ;
      RECT 129.92 128.46 130.52 128.66 ;
      RECT 129.92 129.46 130.52 129.66 ;
      RECT 126.68 129.36 130.12 129.56 ;
      RECT 126.68 131.96 130.12 132.16 ;
      RECT 129.92 131.86 130.52 132.06 ;
      RECT 129.92 132.86 130.52 133.06 ;
      RECT 126.68 132.76 130.12 132.96 ;
      RECT 126.68 135.36 130.12 135.56 ;
      RECT 129.92 135.26 130.52 135.46 ;
      RECT 129.92 136.26 130.52 136.46 ;
      RECT 126.68 136.16 130.12 136.36 ;
      RECT 126.68 138.76 130.12 138.96 ;
      RECT 129.92 138.66 130.52 138.86 ;
      RECT 129.92 139.66 130.52 139.86 ;
      RECT 126.68 139.56 130.12 139.76 ;
      RECT 126.68 142.16 130.12 142.36 ;
      RECT 129.92 142.06 130.52 142.26 ;
      RECT 129.92 143.06 130.52 143.26 ;
      RECT 126.68 142.96 130.12 143.16 ;
      RECT 126.68 145.56 130.12 145.76 ;
      RECT 129.92 145.46 130.52 145.66 ;
      RECT 129.92 146.46 130.52 146.66 ;
      RECT 126.68 146.36 130.12 146.56 ;
      RECT 126.68 148.96 130.12 149.16 ;
      RECT 129.92 148.86 130.52 149.06 ;
      RECT 129.92 149.86 130.52 150.06 ;
      RECT 126.68 149.76 130.12 149.96 ;
      RECT 126.68 152.36 130.12 152.56 ;
      RECT 129.92 152.26 130.52 152.46 ;
      RECT 129.92 153.26 130.52 153.46 ;
      RECT 126.68 153.16 130.12 153.36 ;
      RECT 126.68 155.76 130.12 155.96 ;
      RECT 129.92 155.66 130.52 155.86 ;
      RECT 129.92 156.66 130.52 156.86 ;
      RECT 126.68 156.56 130.12 156.76 ;
      RECT 126.68 159.16 130.12 159.36 ;
      RECT 129.92 159.06 130.52 159.26 ;
      RECT 129.92 160.06 130.52 160.26 ;
      RECT 126.68 159.96 130.12 160.16 ;
      RECT 126.68 162.56 130.12 162.76 ;
      RECT 129.92 162.46 130.52 162.66 ;
      RECT 129.92 163.46 130.52 163.66 ;
      RECT 126.68 163.36 130.12 163.56 ;
      RECT 126.68 165.96 130.12 166.16 ;
      RECT 129.92 165.86 130.52 166.06 ;
      RECT 129.92 166.86 130.52 167.06 ;
      RECT 126.68 166.76 130.12 166.96 ;
      RECT 126.68 169.36 130.12 169.56 ;
      RECT 129.92 169.26 130.52 169.46 ;
      RECT 129.92 170.26 130.52 170.46 ;
      RECT 126.68 170.16 130.12 170.36 ;
      RECT 126.68 172.76 130.12 172.96 ;
      RECT 129.92 172.66 130.52 172.86 ;
      RECT 129.92 173.66 130.52 173.86 ;
      RECT 126.68 173.56 130.12 173.76 ;
      RECT 126.68 176.16 130.12 176.36 ;
      RECT 129.92 176.06 130.52 176.26 ;
      RECT 129.92 177.06 130.52 177.26 ;
      RECT 126.68 176.96 130.12 177.16 ;
      RECT 126.68 179.56 130.12 179.76 ;
      RECT 129.92 179.46 130.52 179.66 ;
      RECT 129.92 180.46 130.52 180.66 ;
      RECT 126.68 180.36 130.12 180.56 ;
      RECT 126.68 182.96 130.12 183.16 ;
      RECT 129.92 182.86 130.52 183.06 ;
      RECT 129.92 183.86 130.52 184.06 ;
      RECT 126.68 183.76 130.12 183.96 ;
      RECT 126.68 186.36 130.12 186.56 ;
      RECT 129.92 186.26 130.52 186.46 ;
      RECT 129.92 187.26 130.52 187.46 ;
      RECT 126.68 187.16 130.12 187.36 ;
      RECT 126.68 189.76 130.12 189.96 ;
      RECT 129.92 189.66 130.52 189.86 ;
      RECT 129.92 190.66 130.52 190.86 ;
      RECT 126.68 190.56 130.12 190.76 ;
      RECT 126.68 193.16 130.12 193.36 ;
      RECT 129.92 193.06 130.52 193.26 ;
      RECT 129.92 194.06 130.52 194.26 ;
      RECT 126.68 193.96 130.12 194.16 ;
      RECT 126.68 196.56 130.12 196.76 ;
      RECT 129.92 196.46 130.52 196.66 ;
      RECT 129.92 197.46 130.52 197.66 ;
      RECT 126.68 197.36 130.12 197.56 ;
      RECT 126.68 199.96 130.12 200.16 ;
      RECT 129.92 199.86 130.52 200.06 ;
      RECT 129.92 200.86 130.52 201.06 ;
      RECT 126.68 200.76 130.12 200.96 ;
      RECT 126.68 203.36 130.12 203.56 ;
      RECT 129.92 203.26 130.52 203.46 ;
      RECT 129.92 204.26 130.52 204.46 ;
      RECT 126.68 204.16 130.12 204.36 ;
      RECT 126.68 206.76 130.12 206.96 ;
      RECT 129.92 206.66 130.52 206.86 ;
      RECT 129.92 207.66 130.52 207.86 ;
      RECT 126.68 207.56 130.12 207.76 ;
      RECT 126.68 210.16 130.12 210.36 ;
      RECT 129.92 210.06 130.52 210.26 ;
      RECT 129.92 211.06 130.52 211.26 ;
      RECT 126.68 210.96 130.12 211.16 ;
      RECT 126.68 213.56 130.12 213.76 ;
      RECT 129.92 213.46 130.52 213.66 ;
      RECT 129.92 214.46 130.52 214.66 ;
      RECT 126.68 214.36 130.12 214.56 ;
      RECT 126.68 216.96 130.12 217.16 ;
      RECT 129.92 216.86 130.52 217.06 ;
      RECT 129.92 217.86 130.52 218.06 ;
      RECT 126.68 217.76 130.12 217.96 ;
      RECT 126.68 220.36 130.12 220.56 ;
      RECT 129.92 220.26 130.52 220.46 ;
      RECT 129.92 221.26 130.52 221.46 ;
      RECT 126.68 221.16 130.12 221.36 ;
      RECT 126.68 223.76 130.12 223.96 ;
      RECT 129.92 223.66 130.52 223.86 ;
      RECT 129.92 224.66 130.52 224.86 ;
      RECT 126.68 224.56 130.12 224.76 ;
      RECT 126.68 227.16 130.12 227.36 ;
      RECT 129.92 227.06 130.52 227.26 ;
      RECT 129.92 228.06 130.52 228.26 ;
      RECT 126.68 227.96 130.12 228.16 ;
      RECT 126.68 230.56 130.12 230.76 ;
      RECT 129.92 230.46 130.52 230.66 ;
      RECT 129.92 231.46 130.52 231.66 ;
      RECT 126.68 231.36 130.12 231.56 ;
      RECT 126.68 233.96 130.12 234.16 ;
      RECT 129.92 233.86 130.52 234.06 ;
      RECT 129.92 234.86 130.52 235.06 ;
      RECT 126.68 234.76 130.12 234.96 ;
      RECT 126.68 237.36 130.12 237.56 ;
      RECT 129.92 237.26 130.52 237.46 ;
      RECT 129.92 238.26 130.52 238.46 ;
      RECT 126.68 238.16 130.12 238.36 ;
      RECT 126.68 240.76 130.12 240.96 ;
      RECT 129.92 240.66 130.52 240.86 ;
      RECT 129.92 241.66 130.52 241.86 ;
      RECT 126.68 241.56 130.12 241.76 ;
      RECT 126.68 244.16 130.12 244.36 ;
      RECT 129.92 244.06 130.52 244.26 ;
      RECT 129.92 245.06 130.52 245.26 ;
      RECT 126.68 244.96 130.12 245.16 ;
      RECT 126.68 247.56 130.12 247.76 ;
      RECT 129.92 247.46 130.52 247.66 ;
      RECT 129.92 248.46 130.52 248.66 ;
      RECT 126.68 248.36 130.12 248.56 ;
      RECT 126.68 250.96 130.12 251.16 ;
      RECT 129.92 250.86 130.52 251.06 ;
      RECT 129.92 251.86 130.52 252.06 ;
      RECT 126.68 251.76 130.12 251.96 ;
      RECT 126.68 254.36 130.12 254.56 ;
      RECT 129.92 254.26 130.52 254.46 ;
      RECT 129.92 255.26 130.52 255.46 ;
      RECT 126.68 255.16 130.12 255.36 ;
      RECT 126.68 257.76 130.12 257.96 ;
      RECT 129.92 257.66 130.52 257.86 ;
      RECT 129.92 258.66 130.52 258.86 ;
      RECT 126.68 258.56 130.12 258.76 ;
      RECT 126.68 261.16 130.12 261.36 ;
      RECT 129.92 261.06 130.52 261.26 ;
      RECT 129.92 262.06 130.52 262.26 ;
      RECT 126.68 261.96 130.12 262.16 ;
      RECT 126.68 264.56 130.12 264.76 ;
      RECT 129.92 264.46 130.52 264.66 ;
      RECT 129.92 265.46 130.52 265.66 ;
      RECT 126.68 265.36 130.12 265.56 ;
      RECT 126.68 267.96 130.12 268.16 ;
      RECT 129.92 267.86 130.52 268.06 ;
      RECT 129.92 268.86 130.52 269.06 ;
      RECT 126.68 268.76 130.12 268.96 ;
      RECT 126.68 271.36 130.12 271.56 ;
      RECT 129.92 271.26 130.52 271.46 ;
      RECT 129.92 272.26 130.52 272.46 ;
      RECT 126.68 272.16 130.12 272.36 ;
      RECT 126.68 274.76 130.12 274.96 ;
      RECT 129.92 274.66 130.52 274.86 ;
      RECT 129.92 275.66 130.52 275.86 ;
      RECT 126.68 275.56 130.12 275.76 ;
      RECT 126.68 278.16 130.12 278.36 ;
      RECT 129.92 278.06 130.52 278.26 ;
      RECT 129.92 279.06 130.52 279.26 ;
      RECT 126.68 278.96 130.12 279.16 ;
      RECT 126.68 281.56 130.12 281.76 ;
      RECT 129.92 281.46 130.52 281.66 ;
      RECT 129.92 282.46 130.52 282.66 ;
      RECT 126.68 282.36 130.12 282.56 ;
      RECT 126.68 284.96 130.12 285.16 ;
      RECT 129.92 284.86 130.52 285.06 ;
      RECT 129.92 285.86 130.52 286.06 ;
      RECT 126.68 285.76 130.12 285.96 ;
      RECT 126.68 288.36 130.12 288.56 ;
      RECT 129.92 288.26 130.52 288.46 ;
      RECT 129.92 289.26 130.52 289.46 ;
      RECT 126.68 289.16 130.12 289.36 ;
      RECT 126.68 291.76 130.12 291.96 ;
      RECT 129.92 291.66 130.52 291.86 ;
      RECT 129.92 292.66 130.52 292.86 ;
      RECT 126.68 292.56 130.12 292.76 ;
      RECT 126.68 295.16 130.12 295.36 ;
      RECT 129.92 295.06 130.52 295.26 ;
      RECT 129.92 296.06 130.52 296.26 ;
      RECT 126.68 295.96 130.12 296.16 ;
      RECT 126.68 298.56 130.12 298.76 ;
      RECT 129.92 298.46 130.52 298.66 ;
      RECT 129.92 299.46 130.52 299.66 ;
      RECT 126.68 299.36 130.12 299.56 ;
      RECT 126.68 301.96 130.12 302.16 ;
      RECT 129.92 301.86 130.52 302.06 ;
      RECT 129.92 302.86 130.52 303.06 ;
      RECT 126.68 302.76 130.12 302.96 ;
      RECT 126.68 305.36 130.12 305.56 ;
      RECT 129.92 305.26 130.52 305.46 ;
      RECT 129.92 306.26 130.52 306.46 ;
      RECT 126.68 306.16 130.12 306.36 ;
      RECT 126.68 308.76 130.12 308.96 ;
      RECT 129.92 308.66 130.52 308.86 ;
      RECT 129.92 309.66 130.52 309.86 ;
      RECT 126.68 309.56 130.12 309.76 ;
      RECT 126.68 312.16 130.12 312.36 ;
      RECT 129.92 312.06 130.52 312.26 ;
      RECT 129.92 313.06 130.52 313.26 ;
      RECT 126.68 312.96 130.12 313.16 ;
      RECT 126.68 315.56 130.12 315.76 ;
      RECT 129.92 315.46 130.52 315.66 ;
      RECT 129.92 316.46 130.52 316.66 ;
      RECT 126.68 316.36 130.12 316.56 ;
      RECT 126.68 318.96 130.12 319.16 ;
      RECT 129.92 318.86 130.52 319.06 ;
      RECT 129.92 319.86 130.52 320.06 ;
      RECT 126.68 319.76 130.12 319.96 ;
      RECT 126.68 322.36 130.12 322.56 ;
      RECT 129.92 322.26 130.52 322.46 ;
      RECT 129.92 323.26 130.52 323.46 ;
      RECT 126.68 323.16 130.12 323.36 ;
      RECT 126.68 325.76 130.12 325.96 ;
      RECT 129.92 325.66 130.52 325.86 ;
      RECT 129.92 326.66 130.52 326.86 ;
      RECT 126.68 326.56 130.12 326.76 ;
      RECT 126.68 329.16 130.12 329.36 ;
      RECT 129.92 329.06 130.52 329.26 ;
      RECT 129.92 330.06 130.52 330.26 ;
      RECT 126.68 329.96 130.12 330.16 ;
      RECT 126.68 332.56 130.12 332.76 ;
      RECT 129.92 332.46 130.52 332.66 ;
      RECT 129.92 333.46 130.52 333.66 ;
      RECT 126.68 333.36 130.12 333.56 ;
      RECT 126.68 335.96 130.12 336.16 ;
      RECT 129.92 335.86 130.52 336.06 ;
      RECT 129.92 336.86 130.52 337.06 ;
      RECT 126.68 336.76 130.12 336.96 ;
      RECT 126.68 339.36 130.12 339.56 ;
      RECT 129.92 339.26 130.52 339.46 ;
      RECT 129.92 340.26 130.52 340.46 ;
      RECT 126.68 340.16 130.12 340.36 ;
      RECT 126.68 342.76 130.12 342.96 ;
      RECT 129.92 342.66 130.52 342.86 ;
      RECT 129.92 343.66 130.52 343.86 ;
      RECT 126.68 343.56 130.12 343.76 ;
      RECT 126.68 346.16 130.12 346.36 ;
      RECT 129.92 346.06 130.52 346.26 ;
      RECT 129.92 347.06 130.52 347.26 ;
      RECT 126.68 346.96 130.12 347.16 ;
      RECT 126.68 349.56 130.12 349.76 ;
      RECT 129.92 349.46 130.52 349.66 ;
      RECT 129.92 350.46 130.52 350.66 ;
      RECT 126.68 350.36 130.12 350.56 ;
      RECT 126.68 352.96 130.12 353.16 ;
      RECT 129.92 352.86 130.52 353.06 ;
      RECT 129.92 353.86 130.52 354.06 ;
      RECT 126.68 353.76 130.12 353.96 ;
      RECT 126.68 356.36 130.12 356.56 ;
      RECT 129.92 356.26 130.52 356.46 ;
      RECT 129.92 357.26 130.52 357.46 ;
      RECT 126.68 357.16 130.12 357.36 ;
      RECT 126.68 359.76 130.12 359.96 ;
      RECT 129.92 359.66 130.52 359.86 ;
      RECT 129.92 360.66 130.52 360.86 ;
      RECT 126.68 360.56 130.12 360.76 ;
      RECT 126.68 363.16 130.12 363.36 ;
      RECT 129.92 363.06 130.52 363.26 ;
      RECT 129.92 364.06 130.52 364.26 ;
      RECT 126.68 363.96 130.12 364.16 ;
      RECT 126.68 366.56 130.12 366.76 ;
      RECT 129.92 366.46 130.52 366.66 ;
      RECT 129.92 367.46 130.52 367.66 ;
      RECT 126.68 367.36 130.12 367.56 ;
      RECT 126.68 369.96 130.12 370.16 ;
      RECT 129.92 369.86 130.52 370.06 ;
      RECT 129.92 370.86 130.52 371.06 ;
      RECT 126.68 370.76 130.12 370.96 ;
      RECT 126.68 373.36 130.12 373.56 ;
      RECT 129.92 373.26 130.52 373.46 ;
      RECT 129.92 374.26 130.52 374.46 ;
      RECT 126.68 374.16 130.12 374.36 ;
      RECT 126.68 376.76 130.12 376.96 ;
      RECT 129.92 376.66 130.52 376.86 ;
      RECT 129.92 377.66 130.52 377.86 ;
      RECT 126.68 377.56 130.12 377.76 ;
      RECT 126.68 380.16 130.12 380.36 ;
      RECT 129.92 380.06 130.52 380.26 ;
      RECT 129.92 381.06 130.52 381.26 ;
      RECT 126.68 380.96 130.12 381.16 ;
      RECT 126.68 383.56 130.12 383.76 ;
      RECT 129.92 383.46 130.52 383.66 ;
      RECT 129.92 384.46 130.52 384.66 ;
      RECT 126.68 384.36 130.12 384.56 ;
      RECT 126.68 386.96 130.12 387.16 ;
      RECT 129.92 386.86 130.52 387.06 ;
      RECT 129.92 387.86 130.52 388.06 ;
      RECT 126.68 387.76 130.12 387.96 ;
      RECT 126.68 390.36 130.12 390.56 ;
      RECT 129.92 390.26 130.52 390.46 ;
      RECT 129.92 391.26 130.52 391.46 ;
      RECT 126.68 391.16 130.12 391.36 ;
      RECT 126.68 393.76 130.12 393.96 ;
      RECT 129.92 393.66 130.52 393.86 ;
      RECT 129.92 394.66 130.52 394.86 ;
      RECT 126.68 394.56 130.12 394.76 ;
      RECT 126.68 397.16 130.12 397.36 ;
      RECT 129.92 397.06 130.52 397.26 ;
      RECT 129.92 398.06 130.52 398.26 ;
      RECT 126.68 397.96 130.12 398.16 ;
      RECT 126.68 400.56 130.12 400.76 ;
      RECT 129.92 400.46 130.52 400.66 ;
      RECT 129.92 401.46 130.52 401.66 ;
      RECT 126.68 401.36 130.12 401.56 ;
      RECT 126.68 403.96 130.12 404.16 ;
      RECT 129.92 403.86 130.52 404.06 ;
      RECT 129.92 404.86 130.52 405.06 ;
      RECT 126.68 404.76 130.12 404.96 ;
      RECT 126.68 407.36 130.12 407.56 ;
      RECT 129.92 407.26 130.52 407.46 ;
      RECT 129.92 408.26 130.52 408.46 ;
      RECT 126.68 408.16 130.12 408.36 ;
      RECT 126.68 410.76 130.12 410.96 ;
      RECT 129.92 410.66 130.52 410.86 ;
      RECT 129.92 411.66 130.52 411.86 ;
      RECT 126.68 411.56 130.12 411.76 ;
      RECT 126.68 414.16 130.12 414.36 ;
      RECT 129.92 414.06 130.52 414.26 ;
      RECT 129.92 415.06 130.52 415.26 ;
      RECT 126.68 414.96 130.12 415.16 ;
      RECT 126.68 417.56 130.12 417.76 ;
      RECT 129.92 417.46 130.52 417.66 ;
      RECT 129.92 418.46 130.52 418.66 ;
      RECT 126.68 418.36 130.12 418.56 ;
      RECT 126.68 420.96 130.12 421.16 ;
      RECT 129.92 420.86 130.52 421.06 ;
      RECT 129.92 421.86 130.52 422.06 ;
      RECT 126.68 421.76 130.12 421.96 ;
      RECT 126.68 424.36 130.12 424.56 ;
      RECT 129.92 424.26 130.52 424.46 ;
      RECT 129.92 425.26 130.52 425.46 ;
      RECT 126.68 425.16 130.12 425.36 ;
      RECT 126.68 427.76 130.12 427.96 ;
      RECT 129.92 427.66 130.52 427.86 ;
      RECT 129.92 428.66 130.52 428.86 ;
      RECT 126.68 428.56 130.12 428.76 ;
      RECT 126.68 431.16 130.12 431.36 ;
      RECT 129.92 431.06 130.52 431.26 ;
      RECT 129.92 432.06 130.52 432.26 ;
      RECT 126.68 431.96 130.12 432.16 ;
      RECT 126.68 434.56 130.12 434.76 ;
      RECT 129.92 434.46 130.52 434.66 ;
      RECT 129.92 435.46 130.52 435.66 ;
      RECT 126.68 435.36 130.12 435.56 ;
      RECT 126.68 437.96 130.12 438.16 ;
      RECT 129.92 437.86 130.52 438.06 ;
      RECT 129.92 438.86 130.52 439.06 ;
      RECT 126.68 438.76 130.12 438.96 ;
      RECT 126.68 441.36 130.12 441.56 ;
      RECT 129.92 441.26 130.52 441.46 ;
      RECT 129.92 442.26 130.52 442.46 ;
      RECT 126.68 442.16 130.12 442.36 ;
      RECT 126.68 444.76 130.12 444.96 ;
      RECT 129.92 444.66 130.52 444.86 ;
      RECT 129.92 445.66 130.52 445.86 ;
      RECT 126.68 445.56 130.12 445.76 ;
      RECT 126.68 448.16 130.12 448.36 ;
      RECT 129.92 448.06 130.52 448.26 ;
      RECT 129.92 449.06 130.52 449.26 ;
      RECT 126.68 448.96 130.12 449.16 ;
      RECT 126.68 451.56 130.12 451.76 ;
      RECT 129.92 451.46 130.52 451.66 ;
      RECT 129.92 452.46 130.52 452.66 ;
      RECT 126.68 452.36 130.12 452.56 ;
      RECT 126.68 454.96 130.12 455.16 ;
      RECT 129.92 454.86 130.52 455.06 ;
      RECT 129.92 455.86 130.52 456.06 ;
      RECT 126.68 455.76 130.12 455.96 ;
      RECT 126.68 458.36 130.12 458.56 ;
      RECT 129.92 458.26 130.52 458.46 ;
      RECT 129.92 459.26 130.52 459.46 ;
      RECT 126.68 459.16 130.12 459.36 ;
      RECT 126.68 461.76 130.12 461.96 ;
      RECT 129.92 461.66 130.52 461.86 ;
      RECT 129.92 462.66 130.52 462.86 ;
      RECT 126.68 462.56 130.12 462.76 ;
      RECT 126.68 465.16 130.12 465.36 ;
      RECT 129.92 465.06 130.52 465.26 ;
      RECT 129.92 466.06 130.52 466.26 ;
      RECT 126.68 465.96 130.12 466.16 ;
      RECT 126.68 468.56 130.12 468.76 ;
      RECT 129.92 468.46 130.52 468.66 ;
      RECT 129.92 469.46 130.52 469.66 ;
      RECT 126.68 469.36 130.12 469.56 ;
      RECT 126.68 471.96 130.12 472.16 ;
      RECT 129.92 471.86 130.52 472.06 ;
      RECT 129.92 472.86 130.52 473.06 ;
      RECT 126.68 472.76 130.12 472.96 ;
      RECT 126.68 475.36 130.12 475.56 ;
      RECT 129.92 475.26 130.52 475.46 ;
      RECT 129.92 476.26 130.52 476.46 ;
      RECT 126.68 476.16 130.12 476.36 ;
      RECT 126.68 478.76 130.12 478.96 ;
      RECT 129.92 478.66 130.52 478.86 ;
      RECT 129.92 479.66 130.52 479.86 ;
      RECT 126.68 479.56 130.12 479.76 ;
      RECT 126.68 482.16 130.12 482.36 ;
      RECT 129.92 482.06 130.52 482.26 ;
      RECT 129.92 483.06 130.52 483.26 ;
      RECT 126.68 482.96 130.12 483.16 ;
      RECT 126.68 485.56 130.12 485.76 ;
      RECT 129.92 485.46 130.52 485.66 ;
      RECT 129.92 486.46 130.52 486.66 ;
      RECT 126.68 486.36 130.12 486.56 ;
      RECT 126.68 488.96 130.12 489.16 ;
      RECT 129.92 488.86 130.52 489.06 ;
      RECT 129.92 489.86 130.52 490.06 ;
      RECT 126.68 489.76 130.12 489.96 ;
      RECT 126.68 492.36 130.12 492.56 ;
      RECT 129.92 492.26 130.52 492.46 ;
      RECT 129.92 493.26 130.52 493.46 ;
      RECT 126.68 493.16 130.12 493.36 ;
      RECT 126.68 495.76 130.12 495.96 ;
      RECT 129.92 495.66 130.52 495.86 ;
      RECT 129.92 496.66 130.52 496.86 ;
      RECT 126.68 496.56 130.12 496.76 ;
      RECT 126.68 499.16 130.12 499.36 ;
      RECT 129.92 499.06 130.52 499.26 ;
      RECT 129.92 500.06 130.52 500.26 ;
      RECT 126.68 499.96 130.12 500.16 ;
      RECT 126.68 502.56 130.12 502.76 ;
      RECT 129.92 502.46 130.52 502.66 ;
      RECT 129.92 503.46 130.52 503.66 ;
      RECT 126.68 503.36 130.12 503.56 ;
      RECT 128.82 37.14 129.02 38.38 ;
      RECT 123.4 37.14 123.6 38.38 ;
      RECT 123.4 37.14 129.02 37.34 ;
      RECT 122.02 37.18 122.22 38.38 ;
      RECT 116.6 37.18 116.8 38.38 ;
      RECT 116.6 37.18 122.22 37.38 ;
      RECT 110.21 38.64 121.81 38.84 ;
      RECT 121.41 37.58 121.81 38.84 ;
      RECT 117.01 37.58 117.41 38.84 ;
      RECT 114.61 37.58 115.01 38.84 ;
      RECT 110.21 37.58 110.61 38.84 ;
      RECT 109.36 71.36 118.54 71.69 ;
      RECT 117.82 71.21 118.54 71.69 ;
      RECT 117.82 74.23 118.54 74.71 ;
      RECT 109.36 74.23 118.54 74.56 ;
      RECT 109.36 78.16 118.54 78.49 ;
      RECT 117.82 78.01 118.54 78.49 ;
      RECT 117.82 81.03 118.54 81.51 ;
      RECT 109.36 81.03 118.54 81.36 ;
      RECT 109.36 84.96 118.54 85.29 ;
      RECT 117.82 84.81 118.54 85.29 ;
      RECT 117.82 87.83 118.54 88.31 ;
      RECT 109.36 87.83 118.54 88.16 ;
      RECT 109.36 91.76 118.54 92.09 ;
      RECT 117.82 91.61 118.54 92.09 ;
      RECT 117.82 94.63 118.54 95.11 ;
      RECT 109.36 94.63 118.54 94.96 ;
      RECT 109.36 98.56 118.54 98.89 ;
      RECT 117.82 98.41 118.54 98.89 ;
      RECT 117.82 101.43 118.54 101.91 ;
      RECT 109.36 101.43 118.54 101.76 ;
      RECT 109.36 105.36 118.54 105.69 ;
      RECT 117.82 105.21 118.54 105.69 ;
      RECT 117.82 108.23 118.54 108.71 ;
      RECT 109.36 108.23 118.54 108.56 ;
      RECT 109.36 112.16 118.54 112.49 ;
      RECT 117.82 112.01 118.54 112.49 ;
      RECT 117.82 115.03 118.54 115.51 ;
      RECT 109.36 115.03 118.54 115.36 ;
      RECT 109.36 118.96 118.54 119.29 ;
      RECT 117.82 118.81 118.54 119.29 ;
      RECT 117.82 121.83 118.54 122.31 ;
      RECT 109.36 121.83 118.54 122.16 ;
      RECT 109.36 125.76 118.54 126.09 ;
      RECT 117.82 125.61 118.54 126.09 ;
      RECT 117.82 128.63 118.54 129.11 ;
      RECT 109.36 128.63 118.54 128.96 ;
      RECT 109.36 132.56 118.54 132.89 ;
      RECT 117.82 132.41 118.54 132.89 ;
      RECT 117.82 135.43 118.54 135.91 ;
      RECT 109.36 135.43 118.54 135.76 ;
      RECT 109.36 139.36 118.54 139.69 ;
      RECT 117.82 139.21 118.54 139.69 ;
      RECT 117.82 142.23 118.54 142.71 ;
      RECT 109.36 142.23 118.54 142.56 ;
      RECT 109.36 146.16 118.54 146.49 ;
      RECT 117.82 146.01 118.54 146.49 ;
      RECT 117.82 149.03 118.54 149.51 ;
      RECT 109.36 149.03 118.54 149.36 ;
      RECT 109.36 152.96 118.54 153.29 ;
      RECT 117.82 152.81 118.54 153.29 ;
      RECT 117.82 155.83 118.54 156.31 ;
      RECT 109.36 155.83 118.54 156.16 ;
      RECT 109.36 159.76 118.54 160.09 ;
      RECT 117.82 159.61 118.54 160.09 ;
      RECT 117.82 162.63 118.54 163.11 ;
      RECT 109.36 162.63 118.54 162.96 ;
      RECT 109.36 166.56 118.54 166.89 ;
      RECT 117.82 166.41 118.54 166.89 ;
      RECT 117.82 169.43 118.54 169.91 ;
      RECT 109.36 169.43 118.54 169.76 ;
      RECT 109.36 173.36 118.54 173.69 ;
      RECT 117.82 173.21 118.54 173.69 ;
      RECT 117.82 176.23 118.54 176.71 ;
      RECT 109.36 176.23 118.54 176.56 ;
      RECT 109.36 180.16 118.54 180.49 ;
      RECT 117.82 180.01 118.54 180.49 ;
      RECT 117.82 183.03 118.54 183.51 ;
      RECT 109.36 183.03 118.54 183.36 ;
      RECT 109.36 186.96 118.54 187.29 ;
      RECT 117.82 186.81 118.54 187.29 ;
      RECT 117.82 189.83 118.54 190.31 ;
      RECT 109.36 189.83 118.54 190.16 ;
      RECT 109.36 193.76 118.54 194.09 ;
      RECT 117.82 193.61 118.54 194.09 ;
      RECT 117.82 196.63 118.54 197.11 ;
      RECT 109.36 196.63 118.54 196.96 ;
      RECT 109.36 200.56 118.54 200.89 ;
      RECT 117.82 200.41 118.54 200.89 ;
      RECT 117.82 203.43 118.54 203.91 ;
      RECT 109.36 203.43 118.54 203.76 ;
      RECT 109.36 207.36 118.54 207.69 ;
      RECT 117.82 207.21 118.54 207.69 ;
      RECT 117.82 210.23 118.54 210.71 ;
      RECT 109.36 210.23 118.54 210.56 ;
      RECT 109.36 214.16 118.54 214.49 ;
      RECT 117.82 214.01 118.54 214.49 ;
      RECT 117.82 217.03 118.54 217.51 ;
      RECT 109.36 217.03 118.54 217.36 ;
      RECT 109.36 220.96 118.54 221.29 ;
      RECT 117.82 220.81 118.54 221.29 ;
      RECT 117.82 223.83 118.54 224.31 ;
      RECT 109.36 223.83 118.54 224.16 ;
      RECT 109.36 227.76 118.54 228.09 ;
      RECT 117.82 227.61 118.54 228.09 ;
      RECT 117.82 230.63 118.54 231.11 ;
      RECT 109.36 230.63 118.54 230.96 ;
      RECT 109.36 234.56 118.54 234.89 ;
      RECT 117.82 234.41 118.54 234.89 ;
      RECT 117.82 237.43 118.54 237.91 ;
      RECT 109.36 237.43 118.54 237.76 ;
      RECT 109.36 241.36 118.54 241.69 ;
      RECT 117.82 241.21 118.54 241.69 ;
      RECT 117.82 244.23 118.54 244.71 ;
      RECT 109.36 244.23 118.54 244.56 ;
      RECT 109.36 248.16 118.54 248.49 ;
      RECT 117.82 248.01 118.54 248.49 ;
      RECT 117.82 251.03 118.54 251.51 ;
      RECT 109.36 251.03 118.54 251.36 ;
      RECT 109.36 254.96 118.54 255.29 ;
      RECT 117.82 254.81 118.54 255.29 ;
      RECT 117.82 257.83 118.54 258.31 ;
      RECT 109.36 257.83 118.54 258.16 ;
      RECT 109.36 261.76 118.54 262.09 ;
      RECT 117.82 261.61 118.54 262.09 ;
      RECT 117.82 264.63 118.54 265.11 ;
      RECT 109.36 264.63 118.54 264.96 ;
      RECT 109.36 268.56 118.54 268.89 ;
      RECT 117.82 268.41 118.54 268.89 ;
      RECT 117.82 271.43 118.54 271.91 ;
      RECT 109.36 271.43 118.54 271.76 ;
      RECT 109.36 275.36 118.54 275.69 ;
      RECT 117.82 275.21 118.54 275.69 ;
      RECT 117.82 278.23 118.54 278.71 ;
      RECT 109.36 278.23 118.54 278.56 ;
      RECT 109.36 282.16 118.54 282.49 ;
      RECT 117.82 282.01 118.54 282.49 ;
      RECT 117.82 285.03 118.54 285.51 ;
      RECT 109.36 285.03 118.54 285.36 ;
      RECT 109.36 288.96 118.54 289.29 ;
      RECT 117.82 288.81 118.54 289.29 ;
      RECT 117.82 291.83 118.54 292.31 ;
      RECT 109.36 291.83 118.54 292.16 ;
      RECT 109.36 295.76 118.54 296.09 ;
      RECT 117.82 295.61 118.54 296.09 ;
      RECT 117.82 298.63 118.54 299.11 ;
      RECT 109.36 298.63 118.54 298.96 ;
      RECT 109.36 302.56 118.54 302.89 ;
      RECT 117.82 302.41 118.54 302.89 ;
      RECT 117.82 305.43 118.54 305.91 ;
      RECT 109.36 305.43 118.54 305.76 ;
      RECT 109.36 309.36 118.54 309.69 ;
      RECT 117.82 309.21 118.54 309.69 ;
      RECT 117.82 312.23 118.54 312.71 ;
      RECT 109.36 312.23 118.54 312.56 ;
      RECT 109.36 316.16 118.54 316.49 ;
      RECT 117.82 316.01 118.54 316.49 ;
      RECT 117.82 319.03 118.54 319.51 ;
      RECT 109.36 319.03 118.54 319.36 ;
      RECT 109.36 322.96 118.54 323.29 ;
      RECT 117.82 322.81 118.54 323.29 ;
      RECT 117.82 325.83 118.54 326.31 ;
      RECT 109.36 325.83 118.54 326.16 ;
      RECT 109.36 329.76 118.54 330.09 ;
      RECT 117.82 329.61 118.54 330.09 ;
      RECT 117.82 332.63 118.54 333.11 ;
      RECT 109.36 332.63 118.54 332.96 ;
      RECT 109.36 336.56 118.54 336.89 ;
      RECT 117.82 336.41 118.54 336.89 ;
      RECT 117.82 339.43 118.54 339.91 ;
      RECT 109.36 339.43 118.54 339.76 ;
      RECT 109.36 343.36 118.54 343.69 ;
      RECT 117.82 343.21 118.54 343.69 ;
      RECT 117.82 346.23 118.54 346.71 ;
      RECT 109.36 346.23 118.54 346.56 ;
      RECT 109.36 350.16 118.54 350.49 ;
      RECT 117.82 350.01 118.54 350.49 ;
      RECT 117.82 353.03 118.54 353.51 ;
      RECT 109.36 353.03 118.54 353.36 ;
      RECT 109.36 356.96 118.54 357.29 ;
      RECT 117.82 356.81 118.54 357.29 ;
      RECT 117.82 359.83 118.54 360.31 ;
      RECT 109.36 359.83 118.54 360.16 ;
      RECT 109.36 363.76 118.54 364.09 ;
      RECT 117.82 363.61 118.54 364.09 ;
      RECT 117.82 366.63 118.54 367.11 ;
      RECT 109.36 366.63 118.54 366.96 ;
      RECT 109.36 370.56 118.54 370.89 ;
      RECT 117.82 370.41 118.54 370.89 ;
      RECT 117.82 373.43 118.54 373.91 ;
      RECT 109.36 373.43 118.54 373.76 ;
      RECT 109.36 377.36 118.54 377.69 ;
      RECT 117.82 377.21 118.54 377.69 ;
      RECT 117.82 380.23 118.54 380.71 ;
      RECT 109.36 380.23 118.54 380.56 ;
      RECT 109.36 384.16 118.54 384.49 ;
      RECT 117.82 384.01 118.54 384.49 ;
      RECT 117.82 387.03 118.54 387.51 ;
      RECT 109.36 387.03 118.54 387.36 ;
      RECT 109.36 390.96 118.54 391.29 ;
      RECT 117.82 390.81 118.54 391.29 ;
      RECT 117.82 393.83 118.54 394.31 ;
      RECT 109.36 393.83 118.54 394.16 ;
      RECT 109.36 397.76 118.54 398.09 ;
      RECT 117.82 397.61 118.54 398.09 ;
      RECT 117.82 400.63 118.54 401.11 ;
      RECT 109.36 400.63 118.54 400.96 ;
      RECT 109.36 404.56 118.54 404.89 ;
      RECT 117.82 404.41 118.54 404.89 ;
      RECT 117.82 407.43 118.54 407.91 ;
      RECT 109.36 407.43 118.54 407.76 ;
      RECT 109.36 411.36 118.54 411.69 ;
      RECT 117.82 411.21 118.54 411.69 ;
      RECT 117.82 414.23 118.54 414.71 ;
      RECT 109.36 414.23 118.54 414.56 ;
      RECT 109.36 418.16 118.54 418.49 ;
      RECT 117.82 418.01 118.54 418.49 ;
      RECT 117.82 421.03 118.54 421.51 ;
      RECT 109.36 421.03 118.54 421.36 ;
      RECT 109.36 424.96 118.54 425.29 ;
      RECT 117.82 424.81 118.54 425.29 ;
      RECT 117.82 427.83 118.54 428.31 ;
      RECT 109.36 427.83 118.54 428.16 ;
      RECT 109.36 431.76 118.54 432.09 ;
      RECT 117.82 431.61 118.54 432.09 ;
      RECT 117.82 434.63 118.54 435.11 ;
      RECT 109.36 434.63 118.54 434.96 ;
      RECT 109.36 438.56 118.54 438.89 ;
      RECT 117.82 438.41 118.54 438.89 ;
      RECT 117.82 441.43 118.54 441.91 ;
      RECT 109.36 441.43 118.54 441.76 ;
      RECT 109.36 445.36 118.54 445.69 ;
      RECT 117.82 445.21 118.54 445.69 ;
      RECT 117.82 448.23 118.54 448.71 ;
      RECT 109.36 448.23 118.54 448.56 ;
      RECT 109.36 452.16 118.54 452.49 ;
      RECT 117.82 452.01 118.54 452.49 ;
      RECT 117.82 455.03 118.54 455.51 ;
      RECT 109.36 455.03 118.54 455.36 ;
      RECT 109.36 458.96 118.54 459.29 ;
      RECT 117.82 458.81 118.54 459.29 ;
      RECT 117.82 461.83 118.54 462.31 ;
      RECT 109.36 461.83 118.54 462.16 ;
      RECT 109.36 465.76 118.54 466.09 ;
      RECT 117.82 465.61 118.54 466.09 ;
      RECT 117.82 468.63 118.54 469.11 ;
      RECT 109.36 468.63 118.54 468.96 ;
      RECT 109.36 472.56 118.54 472.89 ;
      RECT 117.82 472.41 118.54 472.89 ;
      RECT 117.82 475.43 118.54 475.91 ;
      RECT 109.36 475.43 118.54 475.76 ;
      RECT 109.36 479.36 118.54 479.69 ;
      RECT 117.82 479.21 118.54 479.69 ;
      RECT 117.82 482.23 118.54 482.71 ;
      RECT 109.36 482.23 118.54 482.56 ;
      RECT 109.36 486.16 118.54 486.49 ;
      RECT 117.82 486.01 118.54 486.49 ;
      RECT 117.82 489.03 118.54 489.51 ;
      RECT 109.36 489.03 118.54 489.36 ;
      RECT 109.36 492.96 118.54 493.29 ;
      RECT 117.82 492.81 118.54 493.29 ;
      RECT 117.82 495.83 118.54 496.31 ;
      RECT 109.36 495.83 118.54 496.16 ;
      RECT 109.36 499.76 118.54 500.09 ;
      RECT 117.82 499.61 118.54 500.09 ;
      RECT 117.82 502.63 118.54 503.11 ;
      RECT 109.36 502.63 118.54 502.96 ;
      RECT 115.22 37.18 115.42 38.38 ;
      RECT 109.8 37.18 110 38.38 ;
      RECT 109.8 37.18 115.42 37.38 ;
      RECT 108.42 37.18 108.62 38.38 ;
      RECT 103 37.18 103.2 38.38 ;
      RECT 103 37.18 108.62 37.38 ;
      RECT 96.61 38.64 108.21 38.84 ;
      RECT 107.81 37.58 108.21 38.84 ;
      RECT 103.41 37.58 103.81 38.84 ;
      RECT 101.01 37.58 101.41 38.84 ;
      RECT 96.61 37.58 97.01 38.84 ;
      RECT 104.41 510.34 105.51 510.94 ;
      RECT 105.01 68.43 105.41 510.94 ;
      RECT 102.71 510.34 103.81 510.94 ;
      RECT 102.76 68.83 103.16 510.94 ;
      RECT 101.01 510.34 102.11 510.94 ;
      RECT 101.61 68.43 102.01 510.94 ;
      RECT 101.62 37.18 101.82 38.38 ;
      RECT 96.2 37.18 96.4 38.38 ;
      RECT 96.2 37.18 101.82 37.38 ;
      RECT 99.31 510.34 100.41 510.94 ;
      RECT 99.36 68.83 99.76 510.94 ;
      RECT 97.61 510.34 98.71 510.94 ;
      RECT 98.21 68.43 98.61 510.94 ;
      RECT 95.91 510.34 97.01 510.94 ;
      RECT 95.96 68.83 96.36 510.94 ;
      RECT 94.21 510.34 95.31 510.94 ;
      RECT 94.81 68.43 95.21 510.94 ;
      RECT 89.81 38.58 94.61 38.78 ;
      RECT 94.21 37.58 94.61 38.78 ;
      RECT 89.81 37.58 90.21 38.78 ;
      RECT 93.3 37.18 93.61 38.38 ;
      RECT 90.81 37.18 91.12 38.38 ;
      RECT 90.81 37.18 93.61 37.38 ;
      RECT 92.51 510.34 93.61 510.94 ;
      RECT 92.56 68.83 92.96 510.94 ;
      RECT 90.81 510.34 91.91 510.94 ;
      RECT 91.41 68.43 91.81 510.94 ;
      RECT 89.11 510.34 90.21 510.94 ;
      RECT 89.16 68.83 89.56 510.94 ;
      RECT 87.81 510.34 88.61 510.94 ;
      RECT 87.81 69.23 88.19 510.94 ;
      RECT 87.81 69.23 88.67 69.43 ;
      RECT 86.61 510.34 87.41 510.94 ;
      RECT 85.41 510.34 86.21 510.94 ;
      RECT 85.41 510.34 87.41 510.74 ;
      RECT 86.51 68.83 86.71 510.74 ;
      RECT 87.31 68.83 87.51 510.54 ;
      RECT 85.71 65.96 85.91 510.94 ;
      RECT 86.51 68.83 88.65 69.03 ;
      RECT 87.21 67.73 88.51 68.53 ;
      RECT 87.21 66.93 88.01 68.53 ;
      RECT 8.21 10.98 88.01 11.78 ;
      RECT 6.84 10.98 88.01 11.34 ;
      RECT 86.11 65.25 86.31 505.18 ;
      RECT 85.71 65.25 86.31 65.45 ;
      RECT 85.71 63.99 85.91 65.45 ;
      RECT 85.83 58.57 86.03 59.17 ;
      RECT 84.51 58.57 84.71 59.17 ;
      RECT 84.51 58.57 86.03 58.77 ;
      RECT 85.71 37.91 85.91 38.61 ;
      RECT 85.51 37.91 85.91 38.11 ;
      RECT 66.61 38.81 85.31 39.01 ;
      RECT 85.11 37.61 85.31 39.01 ;
      RECT 82.71 37.61 82.91 39.01 ;
      RECT 80.31 37.61 80.51 39.01 ;
      RECT 77.91 37.61 78.11 39.01 ;
      RECT 75.51 37.61 75.71 39.01 ;
      RECT 73.11 37.61 73.31 39.01 ;
      RECT 70.71 37.61 70.91 39.01 ;
      RECT 68.31 37.61 68.51 39.01 ;
      RECT 84.11 63.99 84.31 505.18 ;
      RECT 84.91 63.99 85.11 65.05 ;
      RECT 84.11 63.99 85.11 64.19 ;
      RECT 84.91 65.25 85.11 505.18 ;
      RECT 84.51 65.25 85.11 65.45 ;
      RECT 84.51 64.39 84.71 65.45 ;
      RECT 83.01 510.34 85.01 510.94 ;
      RECT 84.51 65.96 84.71 510.94 ;
      RECT 84.51 37.91 84.71 38.61 ;
      RECT 84.51 37.91 84.91 38.11 ;
      RECT 83.71 63.99 83.91 505.18 ;
      RECT 82.91 63.99 83.11 65.05 ;
      RECT 82.91 63.99 83.91 64.19 ;
      RECT 83.31 37.91 83.51 38.61 ;
      RECT 83.11 37.91 83.51 38.11 ;
      RECT 83.31 58.57 83.51 59.17 ;
      RECT 81.99 58.57 82.19 59.17 ;
      RECT 81.99 58.57 83.51 58.77 ;
      RECT 82.91 65.25 83.11 505.18 ;
      RECT 82.91 65.25 83.51 65.45 ;
      RECT 83.31 64.39 83.51 65.45 ;
      RECT 81.81 510.34 82.61 510.94 ;
      RECT 80.61 510.34 81.41 510.94 ;
      RECT 80.61 510.34 82.61 510.74 ;
      RECT 80.91 65.96 81.11 510.94 ;
      RECT 82.11 37.91 82.31 38.61 ;
      RECT 82.11 37.91 82.51 38.11 ;
      RECT 81.71 65.25 81.91 505.18 ;
      RECT 81.71 65.25 82.31 65.45 ;
      RECT 82.11 63.99 82.31 65.45 ;
      RECT 81.31 65.25 81.51 505.18 ;
      RECT 80.91 65.25 81.51 65.45 ;
      RECT 80.91 63.99 81.11 65.45 ;
      RECT 81.03 58.57 81.23 59.17 ;
      RECT 79.71 58.57 79.91 59.17 ;
      RECT 79.71 58.57 81.23 58.77 ;
      RECT 80.91 37.91 81.11 38.61 ;
      RECT 80.71 37.91 81.11 38.11 ;
      RECT 79.31 63.99 79.51 505.18 ;
      RECT 80.11 63.99 80.31 65.05 ;
      RECT 79.31 63.99 80.31 64.19 ;
      RECT 80.11 65.25 80.31 505.18 ;
      RECT 79.71 65.25 80.31 65.45 ;
      RECT 79.71 64.39 79.91 65.45 ;
      RECT 78.21 510.34 80.21 510.94 ;
      RECT 79.71 65.96 79.91 510.94 ;
      RECT 79.71 37.91 79.91 38.61 ;
      RECT 79.71 37.91 80.11 38.11 ;
      RECT 78.91 63.99 79.11 505.18 ;
      RECT 78.11 63.99 78.31 65.05 ;
      RECT 78.11 63.99 79.11 64.19 ;
      RECT 78.51 37.91 78.71 38.61 ;
      RECT 78.31 37.91 78.71 38.11 ;
      RECT 78.51 58.57 78.71 59.17 ;
      RECT 77.19 58.57 77.39 59.17 ;
      RECT 77.19 58.57 78.71 58.77 ;
      RECT 78.11 65.25 78.31 505.18 ;
      RECT 78.11 65.25 78.71 65.45 ;
      RECT 78.51 64.39 78.71 65.45 ;
      RECT 77.01 510.34 77.81 510.94 ;
      RECT 75.81 510.34 76.61 510.94 ;
      RECT 75.81 510.34 77.81 510.74 ;
      RECT 76.11 65.96 76.31 510.94 ;
      RECT 77.31 37.91 77.51 38.61 ;
      RECT 77.31 37.91 77.71 38.11 ;
      RECT 76.91 65.25 77.11 505.18 ;
      RECT 76.91 65.25 77.51 65.45 ;
      RECT 77.31 63.99 77.51 65.45 ;
      RECT 76.51 65.25 76.71 505.18 ;
      RECT 76.11 65.25 76.71 65.45 ;
      RECT 76.11 63.99 76.31 65.45 ;
      RECT 76.23 58.57 76.43 59.17 ;
      RECT 74.91 58.57 75.11 59.17 ;
      RECT 74.91 58.57 76.43 58.77 ;
      RECT 74.35 24.85 76.41 25.05 ;
      RECT 76.21 24.22 76.41 25.05 ;
      RECT 69.53 12.98 73.21 13.18 ;
      RECT 73.01 12.58 73.21 13.18 ;
      RECT 73.01 12.58 76.31 12.78 ;
      RECT 76.11 37.91 76.31 38.61 ;
      RECT 75.91 37.91 76.31 38.11 ;
      RECT 73.89 23.59 76.27 23.79 ;
      RECT 76.07 22.77 76.27 23.79 ;
      RECT 71.91 22.71 72.11 26.71 ;
      RECT 68.33 22.71 75.69 22.91 ;
      RECT 74.51 63.99 74.71 505.18 ;
      RECT 75.31 63.99 75.51 65.05 ;
      RECT 74.51 63.99 75.51 64.19 ;
      RECT 75.31 65.25 75.51 505.18 ;
      RECT 74.91 65.25 75.51 65.45 ;
      RECT 74.91 64.39 75.11 65.45 ;
      RECT 73.41 510.34 75.41 510.94 ;
      RECT 74.91 65.96 75.11 510.94 ;
      RECT 74.91 37.91 75.11 38.61 ;
      RECT 74.91 37.91 75.31 38.11 ;
      RECT 74.11 63.99 74.31 505.18 ;
      RECT 73.31 63.99 73.51 65.05 ;
      RECT 73.31 63.99 74.31 64.19 ;
      RECT 68.71 16.9 74.28 17.1 ;
      RECT 73.6 15.79 73.8 17.1 ;
      RECT 73.05 15.79 73.8 15.99 ;
      RECT 73.71 37.91 73.91 38.61 ;
      RECT 73.51 37.91 73.91 38.11 ;
      RECT 73.71 58.57 73.91 59.17 ;
      RECT 72.39 58.57 72.59 59.17 ;
      RECT 72.39 58.57 73.91 58.77 ;
      RECT 73.31 65.25 73.51 505.18 ;
      RECT 73.31 65.25 73.91 65.45 ;
      RECT 73.71 64.39 73.91 65.45 ;
      RECT 71.67 16.27 73.4 16.47 ;
      RECT 68.25 16.1 71.87 16.3 ;
      RECT 72.31 23.11 72.51 26.31 ;
      RECT 72.31 23.11 73.11 23.31 ;
      RECT 72.71 26.46 73.11 26.66 ;
      RECT 72.71 24.68 72.91 26.66 ;
      RECT 72.21 510.34 73.01 510.94 ;
      RECT 71.01 510.34 71.81 510.94 ;
      RECT 71.01 510.34 73.01 510.74 ;
      RECT 71.31 65.96 71.51 510.94 ;
      RECT 72.51 37.91 72.71 38.61 ;
      RECT 72.51 37.91 72.91 38.11 ;
      RECT 72.11 65.25 72.31 505.18 ;
      RECT 72.11 65.25 72.71 65.45 ;
      RECT 72.51 63.99 72.71 65.45 ;
      RECT 71.71 65.25 71.91 505.18 ;
      RECT 71.31 65.25 71.91 65.45 ;
      RECT 71.31 63.99 71.51 65.45 ;
      RECT 71.51 23.11 71.71 26.31 ;
      RECT 70.91 23.11 71.71 23.31 ;
      RECT 71.43 58.57 71.63 59.17 ;
      RECT 70.11 58.57 70.31 59.17 ;
      RECT 70.11 58.57 71.63 58.77 ;
      RECT 71.31 37.91 71.51 38.61 ;
      RECT 71.11 37.91 71.51 38.11 ;
      RECT 70.91 26.46 71.31 26.66 ;
      RECT 71.11 24.68 71.31 26.66 ;
      RECT 69.71 63.99 69.91 505.18 ;
      RECT 70.51 63.99 70.71 65.05 ;
      RECT 69.71 63.99 70.71 64.19 ;
      RECT 70.51 65.25 70.71 505.18 ;
      RECT 70.11 65.25 70.71 65.45 ;
      RECT 70.11 64.39 70.31 65.45 ;
      RECT 68.61 510.34 70.61 510.94 ;
      RECT 70.11 65.96 70.31 510.94 ;
      RECT 70.11 37.91 70.31 38.61 ;
      RECT 70.11 37.91 70.51 38.11 ;
      RECT 67.75 23.59 70.13 23.79 ;
      RECT 67.75 22.77 67.95 23.79 ;
      RECT 67.61 24.85 69.67 25.05 ;
      RECT 67.61 24.22 67.81 25.05 ;
      RECT 69.31 63.99 69.51 505.18 ;
      RECT 68.51 63.99 68.71 65.05 ;
      RECT 68.51 63.99 69.51 64.19 ;
      RECT 69.21 15.38 69.41 15.9 ;
      RECT 68.71 15.38 69.41 15.58 ;
      RECT 68.91 37.91 69.11 38.61 ;
      RECT 68.71 37.91 69.11 38.11 ;
      RECT 68.91 58.57 69.11 59.17 ;
      RECT 67.59 58.57 67.79 59.17 ;
      RECT 67.59 58.57 69.11 58.77 ;
      RECT 68.51 65.25 68.71 505.18 ;
      RECT 68.51 65.25 69.11 65.45 ;
      RECT 68.91 64.39 69.11 65.45 ;
      RECT 67.41 510.34 68.21 510.94 ;
      RECT 66.21 510.34 67.01 510.94 ;
      RECT 66.21 510.34 68.21 510.74 ;
      RECT 66.51 65.96 66.71 510.94 ;
      RECT 67.71 37.91 67.91 38.61 ;
      RECT 67.71 37.91 68.11 38.11 ;
      RECT 67.31 65.25 67.51 505.18 ;
      RECT 67.31 65.25 67.91 65.45 ;
      RECT 67.71 63.99 67.91 65.45 ;
      RECT 66.91 65.25 67.11 505.18 ;
      RECT 66.51 65.25 67.11 65.45 ;
      RECT 66.51 63.99 66.71 65.45 ;
      RECT 66.63 58.57 66.83 59.17 ;
      RECT 65.31 58.57 65.51 59.17 ;
      RECT 65.31 58.57 66.83 58.77 ;
      RECT 64.75 24.85 66.81 25.05 ;
      RECT 66.61 24.22 66.81 25.05 ;
      RECT 66.51 37.91 66.71 38.61 ;
      RECT 66.31 37.91 66.71 38.11 ;
      RECT 64.29 23.59 66.67 23.79 ;
      RECT 66.47 22.77 66.67 23.79 ;
      RECT 61.02 16.27 62.75 16.47 ;
      RECT 62.55 16.1 66.17 16.3 ;
      RECT 46.21 38.81 66.11 39.01 ;
      RECT 65.91 37.61 66.11 39.01 ;
      RECT 63.51 37.61 63.71 39.01 ;
      RECT 61.11 37.61 61.31 39.01 ;
      RECT 58.71 37.61 58.91 39.01 ;
      RECT 56.31 37.61 56.51 39.01 ;
      RECT 53.91 37.61 54.11 39.01 ;
      RECT 51.51 37.61 51.71 39.01 ;
      RECT 49.11 37.61 49.31 39.01 ;
      RECT 62.31 22.71 62.51 26.71 ;
      RECT 58.73 22.71 66.09 22.91 ;
      RECT 64.91 63.99 65.11 505.18 ;
      RECT 65.71 63.99 65.91 65.05 ;
      RECT 64.91 63.99 65.91 64.19 ;
      RECT 65.71 65.25 65.91 505.18 ;
      RECT 65.31 65.25 65.91 65.45 ;
      RECT 65.31 64.39 65.51 65.45 ;
      RECT 63.81 510.34 65.81 510.94 ;
      RECT 65.31 65.96 65.51 510.94 ;
      RECT 65.01 15.38 65.21 15.9 ;
      RECT 65.01 15.38 65.71 15.58 ;
      RECT 60.14 16.9 65.71 17.1 ;
      RECT 60.62 15.79 60.82 17.1 ;
      RECT 60.62 15.79 61.37 15.99 ;
      RECT 65.31 37.91 65.51 38.61 ;
      RECT 65.31 37.91 65.71 38.11 ;
      RECT 61.21 12.98 64.89 13.18 ;
      RECT 61.21 12.58 61.41 13.18 ;
      RECT 58.11 12.58 61.41 12.78 ;
      RECT 64.51 63.99 64.71 505.18 ;
      RECT 63.71 63.99 63.91 65.05 ;
      RECT 63.71 63.99 64.71 64.19 ;
      RECT 64.11 37.91 64.31 38.61 ;
      RECT 63.91 37.91 64.31 38.11 ;
      RECT 64.11 58.57 64.31 59.17 ;
      RECT 62.79 58.57 62.99 59.17 ;
      RECT 62.79 58.57 64.31 58.77 ;
      RECT 63.71 65.25 63.91 505.18 ;
      RECT 63.71 65.25 64.31 65.45 ;
      RECT 64.11 64.39 64.31 65.45 ;
      RECT 62.71 23.11 62.91 26.31 ;
      RECT 62.71 23.11 63.51 23.31 ;
      RECT 63.11 26.46 63.51 26.66 ;
      RECT 63.11 24.68 63.31 26.66 ;
      RECT 62.61 510.34 63.41 510.94 ;
      RECT 61.41 510.34 62.21 510.94 ;
      RECT 61.41 510.34 63.41 510.74 ;
      RECT 61.71 65.96 61.91 510.94 ;
      RECT 62.91 37.91 63.11 38.61 ;
      RECT 62.91 37.91 63.31 38.11 ;
      RECT 62.51 65.25 62.71 505.18 ;
      RECT 62.51 65.25 63.11 65.45 ;
      RECT 62.91 63.99 63.11 65.45 ;
      RECT 62.11 65.25 62.31 505.18 ;
      RECT 61.71 65.25 62.31 65.45 ;
      RECT 61.71 63.99 61.91 65.45 ;
      RECT 61.91 23.11 62.11 26.31 ;
      RECT 61.31 23.11 62.11 23.31 ;
      RECT 61.83 58.57 62.03 59.17 ;
      RECT 60.51 58.57 60.71 59.17 ;
      RECT 60.51 58.57 62.03 58.77 ;
      RECT 61.71 37.91 61.91 38.61 ;
      RECT 61.51 37.91 61.91 38.11 ;
      RECT 61.31 26.46 61.71 26.66 ;
      RECT 61.51 24.68 61.71 26.66 ;
      RECT 60.11 63.99 60.31 505.18 ;
      RECT 60.91 63.99 61.11 65.05 ;
      RECT 60.11 63.99 61.11 64.19 ;
      RECT 60.91 65.25 61.11 505.18 ;
      RECT 60.51 65.25 61.11 65.45 ;
      RECT 60.51 64.39 60.71 65.45 ;
      RECT 59.01 510.34 61.01 510.94 ;
      RECT 60.51 65.96 60.71 510.94 ;
      RECT 60.51 37.91 60.71 38.61 ;
      RECT 60.51 37.91 60.91 38.11 ;
      RECT 58.15 23.59 60.53 23.79 ;
      RECT 58.15 22.77 58.35 23.79 ;
      RECT 58.01 24.85 60.07 25.05 ;
      RECT 58.01 24.22 58.21 25.05 ;
      RECT 59.71 63.99 59.91 505.18 ;
      RECT 58.91 63.99 59.11 65.05 ;
      RECT 58.91 63.99 59.91 64.19 ;
      RECT 59.31 37.91 59.51 38.61 ;
      RECT 59.11 37.91 59.51 38.11 ;
      RECT 59.31 58.57 59.51 59.17 ;
      RECT 57.99 58.57 58.19 59.17 ;
      RECT 57.99 58.57 59.51 58.77 ;
      RECT 58.91 65.25 59.11 505.18 ;
      RECT 58.91 65.25 59.51 65.45 ;
      RECT 59.31 64.39 59.51 65.45 ;
      RECT 57.81 510.34 58.61 510.94 ;
      RECT 56.61 510.34 57.41 510.94 ;
      RECT 56.61 510.34 58.61 510.74 ;
      RECT 56.91 65.96 57.11 510.94 ;
      RECT 58.11 37.91 58.31 38.61 ;
      RECT 58.11 37.91 58.51 38.11 ;
      RECT 57.71 65.25 57.91 505.18 ;
      RECT 57.71 65.25 58.31 65.45 ;
      RECT 58.11 63.99 58.31 65.45 ;
      RECT 57.31 65.25 57.51 505.18 ;
      RECT 56.91 65.25 57.51 65.45 ;
      RECT 56.91 63.99 57.11 65.45 ;
      RECT 57.03 58.57 57.23 59.17 ;
      RECT 55.71 58.57 55.91 59.17 ;
      RECT 55.71 58.57 57.23 58.77 ;
      RECT 56.91 37.91 57.11 38.61 ;
      RECT 56.71 37.91 57.11 38.11 ;
      RECT 55.31 63.99 55.51 505.18 ;
      RECT 56.11 63.99 56.31 65.05 ;
      RECT 55.31 63.99 56.31 64.19 ;
      RECT 56.11 65.25 56.31 505.18 ;
      RECT 55.71 65.25 56.31 65.45 ;
      RECT 55.71 64.39 55.91 65.45 ;
      RECT 54.21 510.34 56.21 510.94 ;
      RECT 55.71 65.96 55.91 510.94 ;
      RECT 55.71 37.91 55.91 38.61 ;
      RECT 55.71 37.91 56.11 38.11 ;
      RECT 54.91 63.99 55.11 505.18 ;
      RECT 54.11 63.99 54.31 65.05 ;
      RECT 54.11 63.99 55.11 64.19 ;
      RECT 54.51 37.91 54.71 38.61 ;
      RECT 54.31 37.91 54.71 38.11 ;
      RECT 54.51 58.57 54.71 59.17 ;
      RECT 53.19 58.57 53.39 59.17 ;
      RECT 53.19 58.57 54.71 58.77 ;
      RECT 54.11 65.25 54.31 505.18 ;
      RECT 54.11 65.25 54.71 65.45 ;
      RECT 54.51 64.39 54.71 65.45 ;
      RECT 53.01 510.34 53.81 510.94 ;
      RECT 51.81 510.34 52.61 510.94 ;
      RECT 51.81 510.34 53.81 510.74 ;
      RECT 52.11 65.96 52.31 510.94 ;
      RECT 53.31 37.91 53.51 38.61 ;
      RECT 53.31 37.91 53.71 38.11 ;
      RECT 52.91 65.25 53.11 505.18 ;
      RECT 52.91 65.25 53.51 65.45 ;
      RECT 53.31 63.99 53.51 65.45 ;
      RECT 52.51 65.25 52.71 505.18 ;
      RECT 52.11 65.25 52.71 65.45 ;
      RECT 52.11 63.99 52.31 65.45 ;
      RECT 52.23 58.57 52.43 59.17 ;
      RECT 50.91 58.57 51.11 59.17 ;
      RECT 50.91 58.57 52.43 58.77 ;
      RECT 52.11 37.91 52.31 38.61 ;
      RECT 51.91 37.91 52.31 38.11 ;
      RECT 50.51 63.99 50.71 505.18 ;
      RECT 51.31 63.99 51.51 65.05 ;
      RECT 50.51 63.99 51.51 64.19 ;
      RECT 51.31 65.25 51.51 505.18 ;
      RECT 50.91 65.25 51.51 65.45 ;
      RECT 50.91 64.39 51.11 65.45 ;
      RECT 49.41 510.34 51.41 510.94 ;
      RECT 50.91 65.96 51.11 510.94 ;
      RECT 50.91 37.91 51.11 38.61 ;
      RECT 50.91 37.91 51.31 38.11 ;
      RECT 50.11 63.99 50.31 505.18 ;
      RECT 49.31 63.99 49.51 65.05 ;
      RECT 49.31 63.99 50.31 64.19 ;
      RECT 49.71 37.91 49.91 38.61 ;
      RECT 49.51 37.91 49.91 38.11 ;
      RECT 49.71 58.57 49.91 59.17 ;
      RECT 48.39 58.57 48.59 59.17 ;
      RECT 48.39 58.57 49.91 58.77 ;
      RECT 49.31 65.25 49.51 505.18 ;
      RECT 49.31 65.25 49.91 65.45 ;
      RECT 49.71 64.39 49.91 65.45 ;
      RECT 48.21 510.34 49.01 510.94 ;
      RECT 47.01 510.34 47.81 510.94 ;
      RECT 45.81 510.34 46.61 510.94 ;
      RECT 45.81 510.34 49.01 510.74 ;
      RECT 47.71 68.02 47.91 510.74 ;
      RECT 46.91 68.02 47.11 510.74 ;
      RECT 46.11 65.96 46.31 510.94 ;
      RECT 48.51 37.91 48.71 38.61 ;
      RECT 48.51 37.91 48.91 38.11 ;
      RECT 48.11 65.25 48.31 505.18 ;
      RECT 48.11 65.25 48.71 65.45 ;
      RECT 48.51 63.99 48.71 65.45 ;
      RECT 46.51 65.25 46.71 505.18 ;
      RECT 46.11 65.25 46.71 65.45 ;
      RECT 46.11 63.99 46.31 65.45 ;
      RECT 46.23 58.57 46.43 59.17 ;
      RECT 44.91 58.57 45.11 59.17 ;
      RECT 44.91 58.57 46.43 58.77 ;
      RECT 46.11 37.91 46.31 38.61 ;
      RECT 45.91 37.91 46.31 38.11 ;
      RECT 27.01 38.81 45.71 39.01 ;
      RECT 45.51 37.61 45.71 39.01 ;
      RECT 43.11 37.61 43.31 39.01 ;
      RECT 40.71 37.61 40.91 39.01 ;
      RECT 38.31 37.61 38.51 39.01 ;
      RECT 35.91 37.61 36.11 39.01 ;
      RECT 33.51 37.61 33.71 39.01 ;
      RECT 31.11 37.61 31.31 39.01 ;
      RECT 28.71 37.61 28.91 39.01 ;
      RECT 44.51 63.99 44.71 505.18 ;
      RECT 45.31 63.99 45.51 65.05 ;
      RECT 44.51 63.99 45.51 64.19 ;
      RECT 45.31 65.25 45.51 505.18 ;
      RECT 44.91 65.25 45.51 65.45 ;
      RECT 44.91 64.39 45.11 65.45 ;
      RECT 43.41 510.34 45.41 510.94 ;
      RECT 44.91 65.96 45.11 510.94 ;
      RECT 44.91 37.91 45.11 38.61 ;
      RECT 44.91 37.91 45.31 38.11 ;
      RECT 44.11 63.99 44.31 505.18 ;
      RECT 43.31 63.99 43.51 65.05 ;
      RECT 43.31 63.99 44.31 64.19 ;
      RECT 43.71 37.91 43.91 38.61 ;
      RECT 43.51 37.91 43.91 38.11 ;
      RECT 43.71 58.57 43.91 59.17 ;
      RECT 42.39 58.57 42.59 59.17 ;
      RECT 42.39 58.57 43.91 58.77 ;
      RECT 43.31 65.25 43.51 505.18 ;
      RECT 43.31 65.25 43.91 65.45 ;
      RECT 43.71 64.39 43.91 65.45 ;
      RECT 42.21 510.34 43.01 510.94 ;
      RECT 41.01 510.34 41.81 510.94 ;
      RECT 41.01 510.34 43.01 510.74 ;
      RECT 41.31 65.96 41.51 510.94 ;
      RECT 42.51 37.91 42.71 38.61 ;
      RECT 42.51 37.91 42.91 38.11 ;
      RECT 42.11 65.25 42.31 505.18 ;
      RECT 42.11 65.25 42.71 65.45 ;
      RECT 42.51 63.99 42.71 65.45 ;
      RECT 41.71 65.25 41.91 505.18 ;
      RECT 41.31 65.25 41.91 65.45 ;
      RECT 41.31 63.99 41.51 65.45 ;
      RECT 41.43 58.57 41.63 59.17 ;
      RECT 40.11 58.57 40.31 59.17 ;
      RECT 40.11 58.57 41.63 58.77 ;
      RECT 41.31 37.91 41.51 38.61 ;
      RECT 41.11 37.91 41.51 38.11 ;
      RECT 39.71 63.99 39.91 505.18 ;
      RECT 40.51 63.99 40.71 65.05 ;
      RECT 39.71 63.99 40.71 64.19 ;
      RECT 40.51 65.25 40.71 505.18 ;
      RECT 40.11 65.25 40.71 65.45 ;
      RECT 40.11 64.39 40.31 65.45 ;
      RECT 38.61 510.34 40.61 510.94 ;
      RECT 40.11 65.96 40.31 510.94 ;
      RECT 40.11 37.91 40.31 38.61 ;
      RECT 40.11 37.91 40.51 38.11 ;
      RECT 39.31 63.99 39.51 505.18 ;
      RECT 38.51 63.99 38.71 65.05 ;
      RECT 38.51 63.99 39.51 64.19 ;
      RECT 38.91 37.91 39.11 38.61 ;
      RECT 38.71 37.91 39.11 38.11 ;
      RECT 38.91 58.57 39.11 59.17 ;
      RECT 37.59 58.57 37.79 59.17 ;
      RECT 37.59 58.57 39.11 58.77 ;
      RECT 38.51 65.25 38.71 505.18 ;
      RECT 38.51 65.25 39.11 65.45 ;
      RECT 38.91 64.39 39.11 65.45 ;
      RECT 37.41 510.34 38.21 510.94 ;
      RECT 36.21 510.34 37.01 510.94 ;
      RECT 36.21 510.34 38.21 510.74 ;
      RECT 36.51 65.96 36.71 510.94 ;
      RECT 37.71 37.91 37.91 38.61 ;
      RECT 37.71 37.91 38.11 38.11 ;
      RECT 37.31 65.25 37.51 505.18 ;
      RECT 37.31 65.25 37.91 65.45 ;
      RECT 37.71 63.99 37.91 65.45 ;
      RECT 36.91 65.25 37.11 505.18 ;
      RECT 36.51 65.25 37.11 65.45 ;
      RECT 36.51 63.99 36.71 65.45 ;
      RECT 36.63 58.57 36.83 59.17 ;
      RECT 35.31 58.57 35.51 59.17 ;
      RECT 35.31 58.57 36.83 58.77 ;
      RECT 34.75 24.85 36.81 25.05 ;
      RECT 36.61 24.22 36.81 25.05 ;
      RECT 29.93 12.98 33.61 13.18 ;
      RECT 33.41 12.58 33.61 13.18 ;
      RECT 33.41 12.58 36.71 12.78 ;
      RECT 36.51 37.91 36.71 38.61 ;
      RECT 36.31 37.91 36.71 38.11 ;
      RECT 34.29 23.59 36.67 23.79 ;
      RECT 36.47 22.77 36.67 23.79 ;
      RECT 32.31 22.71 32.51 26.71 ;
      RECT 28.73 22.71 36.09 22.91 ;
      RECT 34.91 63.99 35.11 505.18 ;
      RECT 35.71 63.99 35.91 65.05 ;
      RECT 34.91 63.99 35.91 64.19 ;
      RECT 35.71 65.25 35.91 505.18 ;
      RECT 35.31 65.25 35.91 65.45 ;
      RECT 35.31 64.39 35.51 65.45 ;
      RECT 33.81 510.34 35.81 510.94 ;
      RECT 35.31 65.96 35.51 510.94 ;
      RECT 35.31 37.91 35.51 38.61 ;
      RECT 35.31 37.91 35.71 38.11 ;
      RECT 34.51 63.99 34.71 505.18 ;
      RECT 33.71 63.99 33.91 65.05 ;
      RECT 33.71 63.99 34.71 64.19 ;
      RECT 29.11 16.9 34.68 17.1 ;
      RECT 34 15.79 34.2 17.1 ;
      RECT 33.45 15.79 34.2 15.99 ;
      RECT 34.11 37.91 34.31 38.61 ;
      RECT 33.91 37.91 34.31 38.11 ;
      RECT 34.11 58.57 34.31 59.17 ;
      RECT 32.79 58.57 32.99 59.17 ;
      RECT 32.79 58.57 34.31 58.77 ;
      RECT 33.71 65.25 33.91 505.18 ;
      RECT 33.71 65.25 34.31 65.45 ;
      RECT 34.11 64.39 34.31 65.45 ;
      RECT 32.07 16.27 33.8 16.47 ;
      RECT 28.65 16.1 32.27 16.3 ;
      RECT 32.71 23.11 32.91 26.31 ;
      RECT 32.71 23.11 33.51 23.31 ;
      RECT 33.11 26.46 33.51 26.66 ;
      RECT 33.11 24.68 33.31 26.66 ;
      RECT 32.61 510.34 33.41 510.94 ;
      RECT 31.41 510.34 32.21 510.94 ;
      RECT 31.41 510.34 33.41 510.74 ;
      RECT 31.71 65.96 31.91 510.94 ;
      RECT 32.91 37.91 33.11 38.61 ;
      RECT 32.91 37.91 33.31 38.11 ;
      RECT 32.51 65.25 32.71 505.18 ;
      RECT 32.51 65.25 33.11 65.45 ;
      RECT 32.91 63.99 33.11 65.45 ;
      RECT 32.11 65.25 32.31 505.18 ;
      RECT 31.71 65.25 32.31 65.45 ;
      RECT 31.71 63.99 31.91 65.45 ;
      RECT 31.91 23.11 32.11 26.31 ;
      RECT 31.31 23.11 32.11 23.31 ;
      RECT 31.83 58.57 32.03 59.17 ;
      RECT 30.51 58.57 30.71 59.17 ;
      RECT 30.51 58.57 32.03 58.77 ;
      RECT 31.71 37.91 31.91 38.61 ;
      RECT 31.51 37.91 31.91 38.11 ;
      RECT 31.31 26.46 31.71 26.66 ;
      RECT 31.51 24.68 31.71 26.66 ;
      RECT 30.11 63.99 30.31 505.18 ;
      RECT 30.91 63.99 31.11 65.05 ;
      RECT 30.11 63.99 31.11 64.19 ;
      RECT 30.91 65.25 31.11 505.18 ;
      RECT 30.51 65.25 31.11 65.45 ;
      RECT 30.51 64.39 30.71 65.45 ;
      RECT 29.01 510.34 31.01 510.94 ;
      RECT 30.51 65.96 30.71 510.94 ;
      RECT 30.51 37.91 30.71 38.61 ;
      RECT 30.51 37.91 30.91 38.11 ;
      RECT 28.15 23.59 30.53 23.79 ;
      RECT 28.15 22.77 28.35 23.79 ;
      RECT 28.01 24.85 30.07 25.05 ;
      RECT 28.01 24.22 28.21 25.05 ;
      RECT 29.71 63.99 29.91 505.18 ;
      RECT 28.91 63.99 29.11 65.05 ;
      RECT 28.91 63.99 29.91 64.19 ;
      RECT 29.61 15.38 29.81 15.9 ;
      RECT 29.11 15.38 29.81 15.58 ;
      RECT 29.31 37.91 29.51 38.61 ;
      RECT 29.11 37.91 29.51 38.11 ;
      RECT 29.31 58.57 29.51 59.17 ;
      RECT 27.99 58.57 28.19 59.17 ;
      RECT 27.99 58.57 29.51 58.77 ;
      RECT 28.91 65.25 29.11 505.18 ;
      RECT 28.91 65.25 29.51 65.45 ;
      RECT 29.31 64.39 29.51 65.45 ;
      RECT 27.81 510.34 28.61 510.94 ;
      RECT 26.61 510.34 27.41 510.94 ;
      RECT 26.61 510.34 28.61 510.74 ;
      RECT 26.91 65.96 27.11 510.94 ;
      RECT 28.11 37.91 28.31 38.61 ;
      RECT 28.11 37.91 28.51 38.11 ;
      RECT 27.71 65.25 27.91 505.18 ;
      RECT 27.71 65.25 28.31 65.45 ;
      RECT 28.11 63.99 28.31 65.45 ;
      RECT 27.31 65.25 27.51 505.18 ;
      RECT 26.91 65.25 27.51 65.45 ;
      RECT 26.91 63.99 27.11 65.45 ;
      RECT 27.03 58.57 27.23 59.17 ;
      RECT 25.71 58.57 25.91 59.17 ;
      RECT 25.71 58.57 27.23 58.77 ;
      RECT 25.15 24.85 27.21 25.05 ;
      RECT 27.01 24.22 27.21 25.05 ;
      RECT 26.91 37.91 27.11 38.61 ;
      RECT 26.71 37.91 27.11 38.11 ;
      RECT 24.69 23.59 27.07 23.79 ;
      RECT 26.87 22.77 27.07 23.79 ;
      RECT 21.42 16.27 23.15 16.47 ;
      RECT 22.95 16.1 26.57 16.3 ;
      RECT 7.81 38.81 26.51 39.01 ;
      RECT 26.31 37.61 26.51 39.01 ;
      RECT 23.91 37.61 24.11 39.01 ;
      RECT 21.51 37.61 21.71 39.01 ;
      RECT 19.11 37.61 19.31 39.01 ;
      RECT 16.71 37.61 16.91 39.01 ;
      RECT 14.31 37.61 14.51 39.01 ;
      RECT 11.91 37.61 12.11 39.01 ;
      RECT 9.51 37.61 9.71 39.01 ;
      RECT 22.71 22.71 22.91 26.71 ;
      RECT 19.13 22.71 26.49 22.91 ;
      RECT 25.31 63.99 25.51 505.18 ;
      RECT 26.11 63.99 26.31 65.05 ;
      RECT 25.31 63.99 26.31 64.19 ;
      RECT 26.11 65.25 26.31 505.18 ;
      RECT 25.71 65.25 26.31 65.45 ;
      RECT 25.71 64.39 25.91 65.45 ;
      RECT 24.21 510.34 26.21 510.94 ;
      RECT 25.71 65.96 25.91 510.94 ;
      RECT 25.41 15.38 25.61 15.9 ;
      RECT 25.41 15.38 26.11 15.58 ;
      RECT 20.54 16.9 26.11 17.1 ;
      RECT 21.02 15.79 21.22 17.1 ;
      RECT 21.02 15.79 21.77 15.99 ;
      RECT 25.71 37.91 25.91 38.61 ;
      RECT 25.71 37.91 26.11 38.11 ;
      RECT 21.61 12.98 25.29 13.18 ;
      RECT 21.61 12.58 21.81 13.18 ;
      RECT 18.51 12.58 21.81 12.78 ;
      RECT 24.91 63.99 25.11 505.18 ;
      RECT 24.11 63.99 24.31 65.05 ;
      RECT 24.11 63.99 25.11 64.19 ;
      RECT 24.51 37.91 24.71 38.61 ;
      RECT 24.31 37.91 24.71 38.11 ;
      RECT 24.51 58.57 24.71 59.17 ;
      RECT 23.19 58.57 23.39 59.17 ;
      RECT 23.19 58.57 24.71 58.77 ;
      RECT 24.11 65.25 24.31 505.18 ;
      RECT 24.11 65.25 24.71 65.45 ;
      RECT 24.51 64.39 24.71 65.45 ;
      RECT 23.11 23.11 23.31 26.31 ;
      RECT 23.11 23.11 23.91 23.31 ;
      RECT 23.51 26.46 23.91 26.66 ;
      RECT 23.51 24.68 23.71 26.66 ;
      RECT 23.01 510.34 23.81 510.94 ;
      RECT 21.81 510.34 22.61 510.94 ;
      RECT 21.81 510.34 23.81 510.74 ;
      RECT 22.11 65.96 22.31 510.94 ;
      RECT 23.31 37.91 23.51 38.61 ;
      RECT 23.31 37.91 23.71 38.11 ;
      RECT 22.91 65.25 23.11 505.18 ;
      RECT 22.91 65.25 23.51 65.45 ;
      RECT 23.31 63.99 23.51 65.45 ;
      RECT 22.51 65.25 22.71 505.18 ;
      RECT 22.11 65.25 22.71 65.45 ;
      RECT 22.11 63.99 22.31 65.45 ;
      RECT 22.31 23.11 22.51 26.31 ;
      RECT 21.71 23.11 22.51 23.31 ;
      RECT 22.23 58.57 22.43 59.17 ;
      RECT 20.91 58.57 21.11 59.17 ;
      RECT 20.91 58.57 22.43 58.77 ;
      RECT 22.11 37.91 22.31 38.61 ;
      RECT 21.91 37.91 22.31 38.11 ;
      RECT 21.71 26.46 22.11 26.66 ;
      RECT 21.91 24.68 22.11 26.66 ;
      RECT 20.51 63.99 20.71 505.18 ;
      RECT 21.31 63.99 21.51 65.05 ;
      RECT 20.51 63.99 21.51 64.19 ;
      RECT 21.31 65.25 21.51 505.18 ;
      RECT 20.91 65.25 21.51 65.45 ;
      RECT 20.91 64.39 21.11 65.45 ;
      RECT 19.41 510.34 21.41 510.94 ;
      RECT 20.91 65.96 21.11 510.94 ;
      RECT 20.91 37.91 21.11 38.61 ;
      RECT 20.91 37.91 21.31 38.11 ;
      RECT 18.55 23.59 20.93 23.79 ;
      RECT 18.55 22.77 18.75 23.79 ;
      RECT 18.41 24.85 20.47 25.05 ;
      RECT 18.41 24.22 18.61 25.05 ;
      RECT 20.11 63.99 20.31 505.18 ;
      RECT 19.31 63.99 19.51 65.05 ;
      RECT 19.31 63.99 20.31 64.19 ;
      RECT 19.71 37.91 19.91 38.61 ;
      RECT 19.51 37.91 19.91 38.11 ;
      RECT 19.71 58.57 19.91 59.17 ;
      RECT 18.39 58.57 18.59 59.17 ;
      RECT 18.39 58.57 19.91 58.77 ;
      RECT 19.31 65.25 19.51 505.18 ;
      RECT 19.31 65.25 19.91 65.45 ;
      RECT 19.71 64.39 19.91 65.45 ;
      RECT 18.21 510.34 19.01 510.94 ;
      RECT 17.01 510.34 17.81 510.94 ;
      RECT 17.01 510.34 19.01 510.74 ;
      RECT 17.31 65.96 17.51 510.94 ;
      RECT 18.51 37.91 18.71 38.61 ;
      RECT 18.51 37.91 18.91 38.11 ;
      RECT 18.11 65.25 18.31 505.18 ;
      RECT 18.11 65.25 18.71 65.45 ;
      RECT 18.51 63.99 18.71 65.45 ;
      RECT 17.71 65.25 17.91 505.18 ;
      RECT 17.31 65.25 17.91 65.45 ;
      RECT 17.31 63.99 17.51 65.45 ;
      RECT 17.43 58.57 17.63 59.17 ;
      RECT 16.11 58.57 16.31 59.17 ;
      RECT 16.11 58.57 17.63 58.77 ;
      RECT 17.31 37.91 17.51 38.61 ;
      RECT 17.11 37.91 17.51 38.11 ;
      RECT 15.71 63.99 15.91 505.18 ;
      RECT 16.51 63.99 16.71 65.05 ;
      RECT 15.71 63.99 16.71 64.19 ;
      RECT 16.51 65.25 16.71 505.18 ;
      RECT 16.11 65.25 16.71 65.45 ;
      RECT 16.11 64.39 16.31 65.45 ;
      RECT 14.61 510.34 16.61 510.94 ;
      RECT 16.11 65.96 16.31 510.94 ;
      RECT 16.11 37.91 16.31 38.61 ;
      RECT 16.11 37.91 16.51 38.11 ;
      RECT 15.31 63.99 15.51 505.18 ;
      RECT 14.51 63.99 14.71 65.05 ;
      RECT 14.51 63.99 15.51 64.19 ;
      RECT 14.91 37.91 15.11 38.61 ;
      RECT 14.71 37.91 15.11 38.11 ;
      RECT 14.91 58.57 15.11 59.17 ;
      RECT 13.59 58.57 13.79 59.17 ;
      RECT 13.59 58.57 15.11 58.77 ;
      RECT 14.51 65.25 14.71 505.18 ;
      RECT 14.51 65.25 15.11 65.45 ;
      RECT 14.91 64.39 15.11 65.45 ;
      RECT 13.41 510.34 14.21 510.94 ;
      RECT 12.21 510.34 13.01 510.94 ;
      RECT 12.21 510.34 14.21 510.74 ;
      RECT 12.51 65.96 12.71 510.94 ;
      RECT 13.71 37.91 13.91 38.61 ;
      RECT 13.71 37.91 14.11 38.11 ;
      RECT 13.31 65.25 13.51 505.18 ;
      RECT 13.31 65.25 13.91 65.45 ;
      RECT 13.71 63.99 13.91 65.45 ;
      RECT 12.91 65.25 13.11 505.18 ;
      RECT 12.51 65.25 13.11 65.45 ;
      RECT 12.51 63.99 12.71 65.45 ;
      RECT 12.63 58.57 12.83 59.17 ;
      RECT 11.31 58.57 11.51 59.17 ;
      RECT 11.31 58.57 12.83 58.77 ;
      RECT 12.51 37.91 12.71 38.61 ;
      RECT 12.31 37.91 12.71 38.11 ;
      RECT 10.91 63.99 11.11 505.18 ;
      RECT 11.71 63.99 11.91 65.05 ;
      RECT 10.91 63.99 11.91 64.19 ;
      RECT 11.71 65.25 11.91 505.18 ;
      RECT 11.31 65.25 11.91 65.45 ;
      RECT 11.31 64.39 11.51 65.45 ;
      RECT 9.81 510.34 11.81 510.94 ;
      RECT 11.31 65.96 11.51 510.94 ;
      RECT 11.31 37.91 11.51 38.61 ;
      RECT 11.31 37.91 11.71 38.11 ;
      RECT 10.51 63.99 10.71 505.18 ;
      RECT 9.71 63.99 9.91 65.05 ;
      RECT 9.71 63.99 10.71 64.19 ;
      RECT 10.11 37.91 10.31 38.61 ;
      RECT 9.91 37.91 10.31 38.11 ;
      RECT 10.11 58.57 10.31 59.17 ;
      RECT 8.79 58.57 8.99 59.17 ;
      RECT 8.79 58.57 10.31 58.77 ;
      RECT 9.71 65.25 9.91 505.18 ;
      RECT 9.71 65.25 10.31 65.45 ;
      RECT 10.11 64.39 10.31 65.45 ;
      RECT 8.61 510.34 9.41 510.94 ;
      RECT 7.41 510.34 8.21 510.94 ;
      RECT 7.21 510.34 9.41 510.74 ;
      RECT 8.11 68.04 8.31 510.74 ;
      RECT 7.31 68.04 7.51 510.74 ;
      RECT 6.24 506.6 7.51 508.6 ;
      RECT 6.24 502.66 7.51 503.46 ;
      RECT 6.24 499.26 7.51 500.06 ;
      RECT 6.24 495.86 7.51 496.66 ;
      RECT 6.24 492.46 7.51 493.26 ;
      RECT 6.24 489.06 7.51 489.86 ;
      RECT 6.24 485.66 7.51 486.46 ;
      RECT 6.24 482.26 7.51 483.06 ;
      RECT 6.24 478.86 7.51 479.66 ;
      RECT 6.24 475.46 7.51 476.26 ;
      RECT 6.24 472.06 7.51 472.86 ;
      RECT 6.24 468.66 7.51 469.46 ;
      RECT 6.24 465.26 7.51 466.06 ;
      RECT 6.24 461.86 7.51 462.66 ;
      RECT 6.24 458.46 7.51 459.26 ;
      RECT 6.24 455.06 7.51 455.86 ;
      RECT 6.24 451.66 7.51 452.46 ;
      RECT 6.24 448.26 7.51 449.06 ;
      RECT 6.24 444.86 7.51 445.66 ;
      RECT 6.24 441.46 7.51 442.26 ;
      RECT 6.24 438.06 7.51 438.86 ;
      RECT 6.24 434.66 7.51 435.46 ;
      RECT 6.24 431.26 7.51 432.06 ;
      RECT 6.24 427.86 7.51 428.66 ;
      RECT 6.24 424.46 7.51 425.26 ;
      RECT 6.24 421.06 7.51 421.86 ;
      RECT 6.24 417.66 7.51 418.46 ;
      RECT 6.24 414.26 7.51 415.06 ;
      RECT 6.24 410.86 7.51 411.66 ;
      RECT 6.24 407.46 7.51 408.26 ;
      RECT 6.24 404.06 7.51 404.86 ;
      RECT 6.24 400.66 7.51 401.46 ;
      RECT 6.24 397.26 7.51 398.06 ;
      RECT 6.24 393.86 7.51 394.66 ;
      RECT 6.24 390.46 7.51 391.26 ;
      RECT 6.24 387.06 7.51 387.86 ;
      RECT 6.24 383.66 7.51 384.46 ;
      RECT 6.24 380.26 7.51 381.06 ;
      RECT 6.24 376.86 7.51 377.66 ;
      RECT 6.24 373.46 7.51 374.26 ;
      RECT 6.24 370.06 7.51 370.86 ;
      RECT 6.24 366.66 7.51 367.46 ;
      RECT 6.24 363.26 7.51 364.06 ;
      RECT 6.24 359.86 7.51 360.66 ;
      RECT 6.24 356.46 7.51 357.26 ;
      RECT 6.24 353.06 7.51 353.86 ;
      RECT 6.24 349.66 7.51 350.46 ;
      RECT 6.24 346.26 7.51 347.06 ;
      RECT 6.24 342.86 7.51 343.66 ;
      RECT 6.24 339.46 7.51 340.26 ;
      RECT 6.24 336.06 7.51 336.86 ;
      RECT 6.24 332.66 7.51 333.46 ;
      RECT 6.24 329.26 7.51 330.06 ;
      RECT 6.24 325.86 7.51 326.66 ;
      RECT 6.24 322.46 7.51 323.26 ;
      RECT 6.24 319.06 7.51 319.86 ;
      RECT 6.24 315.66 7.51 316.46 ;
      RECT 6.24 312.26 7.51 313.06 ;
      RECT 6.24 308.86 7.51 309.66 ;
      RECT 6.24 305.46 7.51 306.26 ;
      RECT 6.24 302.06 7.51 302.86 ;
      RECT 6.24 298.66 7.51 299.46 ;
      RECT 6.24 295.26 7.51 296.06 ;
      RECT 6.24 291.86 7.51 292.66 ;
      RECT 6.24 288.46 7.51 289.26 ;
      RECT 6.24 285.06 7.51 285.86 ;
      RECT 6.24 281.66 7.51 282.46 ;
      RECT 6.24 278.26 7.51 279.06 ;
      RECT 6.24 274.86 7.51 275.66 ;
      RECT 6.24 271.46 7.51 272.26 ;
      RECT 6.24 268.06 7.51 268.86 ;
      RECT 6.24 264.66 7.51 265.46 ;
      RECT 6.24 261.26 7.51 262.06 ;
      RECT 6.24 257.86 7.51 258.66 ;
      RECT 6.24 254.46 7.51 255.26 ;
      RECT 6.24 251.06 7.51 251.86 ;
      RECT 6.24 247.66 7.51 248.46 ;
      RECT 6.24 244.26 7.51 245.06 ;
      RECT 6.24 240.86 7.51 241.66 ;
      RECT 6.24 237.46 7.51 238.26 ;
      RECT 6.24 234.06 7.51 234.86 ;
      RECT 6.24 230.66 7.51 231.46 ;
      RECT 6.24 227.26 7.51 228.06 ;
      RECT 6.24 223.86 7.51 224.66 ;
      RECT 6.24 220.46 7.51 221.26 ;
      RECT 6.24 217.06 7.51 217.86 ;
      RECT 6.24 213.66 7.51 214.46 ;
      RECT 6.24 210.26 7.51 211.06 ;
      RECT 6.24 206.86 7.51 207.66 ;
      RECT 6.24 203.46 7.51 204.26 ;
      RECT 6.24 200.06 7.51 200.86 ;
      RECT 6.24 196.66 7.51 197.46 ;
      RECT 6.24 193.26 7.51 194.06 ;
      RECT 6.24 189.86 7.51 190.66 ;
      RECT 6.24 186.46 7.51 187.26 ;
      RECT 6.24 183.06 7.51 183.86 ;
      RECT 6.24 179.66 7.51 180.46 ;
      RECT 6.24 176.26 7.51 177.06 ;
      RECT 6.24 172.86 7.51 173.66 ;
      RECT 6.24 169.46 7.51 170.26 ;
      RECT 6.24 166.06 7.51 166.86 ;
      RECT 6.24 162.66 7.51 163.46 ;
      RECT 6.24 159.26 7.51 160.06 ;
      RECT 6.24 155.86 7.51 156.66 ;
      RECT 6.24 152.46 7.51 153.26 ;
      RECT 6.24 149.06 7.51 149.86 ;
      RECT 6.24 145.66 7.51 146.46 ;
      RECT 6.24 142.26 7.51 143.06 ;
      RECT 6.24 138.86 7.51 139.66 ;
      RECT 6.24 135.46 7.51 136.26 ;
      RECT 6.24 132.06 7.51 132.86 ;
      RECT 6.24 128.66 7.51 129.46 ;
      RECT 6.24 125.26 7.51 126.06 ;
      RECT 6.24 121.86 7.51 122.66 ;
      RECT 6.24 118.46 7.51 119.26 ;
      RECT 6.24 115.06 7.51 115.86 ;
      RECT 6.24 111.66 7.51 112.46 ;
      RECT 6.24 108.26 7.51 109.06 ;
      RECT 6.24 104.86 7.51 105.66 ;
      RECT 6.24 101.46 7.51 102.26 ;
      RECT 6.24 98.06 7.51 98.86 ;
      RECT 6.24 94.66 7.51 95.46 ;
      RECT 6.24 91.26 7.51 92.06 ;
      RECT 6.24 87.86 7.51 88.66 ;
      RECT 6.24 84.46 7.51 85.26 ;
      RECT 6.24 81.06 7.51 81.86 ;
      RECT 6.24 77.66 7.51 78.46 ;
      RECT 6.24 74.26 7.51 75.06 ;
      RECT 6.24 70.86 7.51 71.66 ;
      RECT 7.31 68.04 8.31 68.24 ;
      RECT 8.91 37.91 9.11 38.61 ;
      RECT 8.91 37.91 9.31 38.11 ;
      RECT 8.51 65.25 8.71 505.18 ;
      RECT 8.51 65.25 9.11 65.45 ;
      RECT 8.91 63.99 9.11 65.45 ;
      RECT 233.76 12.64 234.36 13.74 ;
      RECT 153.45 31.13 234.36 32.13 ;
      RECT 6.24 41.29 234.36 42.29 ;
      RECT 6.24 50.24 234.36 51.24 ;
      RECT 6.24 54.22 234.36 55.22 ;
      RECT 140.89 57.02 234.36 58.02 ;
      RECT 233.76 69.16 234.36 69.96 ;
      RECT 233.76 72.56 234.36 73.36 ;
      RECT 233.76 75.96 234.36 76.76 ;
      RECT 233.76 79.36 234.36 80.16 ;
      RECT 233.76 82.76 234.36 83.56 ;
      RECT 233.76 86.16 234.36 86.96 ;
      RECT 233.76 89.56 234.36 90.36 ;
      RECT 233.76 92.96 234.36 93.76 ;
      RECT 233.76 96.36 234.36 97.16 ;
      RECT 233.76 99.76 234.36 100.56 ;
      RECT 233.76 103.16 234.36 103.96 ;
      RECT 233.76 106.56 234.36 107.36 ;
      RECT 233.76 109.96 234.36 110.76 ;
      RECT 233.76 113.36 234.36 114.16 ;
      RECT 233.76 116.76 234.36 117.56 ;
      RECT 233.76 120.16 234.36 120.96 ;
      RECT 233.76 123.56 234.36 124.36 ;
      RECT 233.76 126.96 234.36 127.76 ;
      RECT 233.76 130.36 234.36 131.16 ;
      RECT 233.76 133.76 234.36 134.56 ;
      RECT 233.76 137.16 234.36 137.96 ;
      RECT 233.76 140.56 234.36 141.36 ;
      RECT 233.76 143.96 234.36 144.76 ;
      RECT 233.76 147.36 234.36 148.16 ;
      RECT 233.76 150.76 234.36 151.56 ;
      RECT 233.76 154.16 234.36 154.96 ;
      RECT 233.76 157.56 234.36 158.36 ;
      RECT 233.76 160.96 234.36 161.76 ;
      RECT 233.76 164.36 234.36 165.16 ;
      RECT 233.76 167.76 234.36 168.56 ;
      RECT 233.76 171.16 234.36 171.96 ;
      RECT 233.76 174.56 234.36 175.36 ;
      RECT 233.76 177.96 234.36 178.76 ;
      RECT 233.76 181.36 234.36 182.16 ;
      RECT 233.76 184.76 234.36 185.56 ;
      RECT 233.76 188.16 234.36 188.96 ;
      RECT 233.76 191.56 234.36 192.36 ;
      RECT 233.76 194.96 234.36 195.76 ;
      RECT 233.76 198.36 234.36 199.16 ;
      RECT 233.76 201.76 234.36 202.56 ;
      RECT 233.76 205.16 234.36 205.96 ;
      RECT 233.76 208.56 234.36 209.36 ;
      RECT 233.76 211.96 234.36 212.76 ;
      RECT 233.76 215.36 234.36 216.16 ;
      RECT 233.76 218.76 234.36 219.56 ;
      RECT 233.76 222.16 234.36 222.96 ;
      RECT 233.76 225.56 234.36 226.36 ;
      RECT 233.76 228.96 234.36 229.76 ;
      RECT 233.76 232.36 234.36 233.16 ;
      RECT 233.76 235.76 234.36 236.56 ;
      RECT 233.76 239.16 234.36 239.96 ;
      RECT 233.76 242.56 234.36 243.36 ;
      RECT 233.76 245.96 234.36 246.76 ;
      RECT 233.76 249.36 234.36 250.16 ;
      RECT 233.76 252.76 234.36 253.56 ;
      RECT 233.76 256.16 234.36 256.96 ;
      RECT 233.76 259.56 234.36 260.36 ;
      RECT 233.76 262.96 234.36 263.76 ;
      RECT 233.76 266.36 234.36 267.16 ;
      RECT 233.76 269.76 234.36 270.56 ;
      RECT 233.76 273.16 234.36 273.96 ;
      RECT 233.76 276.56 234.36 277.36 ;
      RECT 233.76 279.96 234.36 280.76 ;
      RECT 233.76 283.36 234.36 284.16 ;
      RECT 233.76 286.76 234.36 287.56 ;
      RECT 233.76 290.16 234.36 290.96 ;
      RECT 233.76 293.56 234.36 294.36 ;
      RECT 233.76 296.96 234.36 297.76 ;
      RECT 233.76 300.36 234.36 301.16 ;
      RECT 233.76 303.76 234.36 304.56 ;
      RECT 233.76 307.16 234.36 307.96 ;
      RECT 233.76 310.56 234.36 311.36 ;
      RECT 233.76 313.96 234.36 314.76 ;
      RECT 233.76 317.36 234.36 318.16 ;
      RECT 233.76 320.76 234.36 321.56 ;
      RECT 233.76 324.16 234.36 324.96 ;
      RECT 233.76 327.56 234.36 328.36 ;
      RECT 233.76 330.96 234.36 331.76 ;
      RECT 233.76 334.36 234.36 335.16 ;
      RECT 233.76 337.76 234.36 338.56 ;
      RECT 233.76 341.16 234.36 341.96 ;
      RECT 233.76 344.56 234.36 345.36 ;
      RECT 233.76 347.96 234.36 348.76 ;
      RECT 233.76 351.36 234.36 352.16 ;
      RECT 233.76 354.76 234.36 355.56 ;
      RECT 233.76 358.16 234.36 358.96 ;
      RECT 233.76 361.56 234.36 362.36 ;
      RECT 233.76 364.96 234.36 365.76 ;
      RECT 233.76 368.36 234.36 369.16 ;
      RECT 233.76 371.76 234.36 372.56 ;
      RECT 233.76 375.16 234.36 375.96 ;
      RECT 233.76 378.56 234.36 379.36 ;
      RECT 233.76 381.96 234.36 382.76 ;
      RECT 233.76 385.36 234.36 386.16 ;
      RECT 233.76 388.76 234.36 389.56 ;
      RECT 233.76 392.16 234.36 392.96 ;
      RECT 233.76 395.56 234.36 396.36 ;
      RECT 233.76 398.96 234.36 399.76 ;
      RECT 233.76 402.36 234.36 403.16 ;
      RECT 233.76 405.76 234.36 406.56 ;
      RECT 233.76 409.16 234.36 409.96 ;
      RECT 233.76 412.56 234.36 413.36 ;
      RECT 233.76 415.96 234.36 416.76 ;
      RECT 233.76 419.36 234.36 420.16 ;
      RECT 233.76 422.76 234.36 423.56 ;
      RECT 233.76 426.16 234.36 426.96 ;
      RECT 233.76 429.56 234.36 430.36 ;
      RECT 233.76 432.96 234.36 433.76 ;
      RECT 233.76 436.36 234.36 437.16 ;
      RECT 233.76 439.76 234.36 440.56 ;
      RECT 233.76 443.16 234.36 443.96 ;
      RECT 233.76 446.56 234.36 447.36 ;
      RECT 233.76 449.96 234.36 450.76 ;
      RECT 233.76 453.36 234.36 454.16 ;
      RECT 233.76 456.76 234.36 457.56 ;
      RECT 233.76 460.16 234.36 460.96 ;
      RECT 233.76 463.56 234.36 464.36 ;
      RECT 233.76 466.96 234.36 467.76 ;
      RECT 233.76 470.36 234.36 471.16 ;
      RECT 233.76 473.76 234.36 474.56 ;
      RECT 233.76 477.16 234.36 477.96 ;
      RECT 233.76 480.56 234.36 481.36 ;
      RECT 233.76 483.96 234.36 484.76 ;
      RECT 233.76 487.36 234.36 488.16 ;
      RECT 233.76 490.76 234.36 491.56 ;
      RECT 233.76 494.16 234.36 494.96 ;
      RECT 233.76 497.56 234.36 498.36 ;
      RECT 233.76 500.96 234.36 501.76 ;
      RECT 233.76 504.36 234.36 505.16 ;
      RECT 233.76 505.6 234.36 506 ;
      RECT 233.76 509 234.36 509.8 ;
      RECT 6.82 9.34 233.78 9.54 ;
      RECT 152.09 19.01 233.77 19.81 ;
      RECT 231.19 6.24 233.19 6.84 ;
      RECT 232.69 68.76 232.89 70.2 ;
      RECT 232.69 70.4 232.89 71.16 ;
      RECT 232.69 71.36 232.89 72.12 ;
      RECT 232.69 72.32 232.89 73.6 ;
      RECT 232.69 73.8 232.89 74.56 ;
      RECT 232.69 74.76 232.89 75.52 ;
      RECT 232.69 75.72 232.89 77 ;
      RECT 232.69 77.2 232.89 77.96 ;
      RECT 232.69 78.16 232.89 78.92 ;
      RECT 232.69 79.12 232.89 80.4 ;
      RECT 232.69 80.6 232.89 81.36 ;
      RECT 232.69 81.56 232.89 82.32 ;
      RECT 232.69 82.52 232.89 83.8 ;
      RECT 232.69 84 232.89 84.76 ;
      RECT 232.69 84.96 232.89 85.72 ;
      RECT 232.69 85.92 232.89 87.2 ;
      RECT 232.69 87.4 232.89 88.16 ;
      RECT 232.69 88.36 232.89 89.12 ;
      RECT 232.69 89.32 232.89 90.6 ;
      RECT 232.69 90.8 232.89 91.56 ;
      RECT 232.69 91.76 232.89 92.52 ;
      RECT 232.69 92.72 232.89 94 ;
      RECT 232.69 94.2 232.89 94.96 ;
      RECT 232.69 95.16 232.89 95.92 ;
      RECT 232.69 96.12 232.89 97.4 ;
      RECT 232.69 97.6 232.89 98.36 ;
      RECT 232.69 98.56 232.89 99.32 ;
      RECT 232.69 99.52 232.89 100.8 ;
      RECT 232.69 101 232.89 101.76 ;
      RECT 232.69 101.96 232.89 102.72 ;
      RECT 232.69 102.92 232.89 104.2 ;
      RECT 232.69 104.4 232.89 105.16 ;
      RECT 232.69 105.36 232.89 106.12 ;
      RECT 232.69 106.32 232.89 107.6 ;
      RECT 232.69 107.8 232.89 108.56 ;
      RECT 232.69 108.76 232.89 109.52 ;
      RECT 232.69 109.72 232.89 111 ;
      RECT 232.69 111.2 232.89 111.96 ;
      RECT 232.69 112.16 232.89 112.92 ;
      RECT 232.69 113.12 232.89 114.4 ;
      RECT 232.69 114.6 232.89 115.36 ;
      RECT 232.69 115.56 232.89 116.32 ;
      RECT 232.69 116.52 232.89 117.8 ;
      RECT 232.69 118 232.89 118.76 ;
      RECT 232.69 118.96 232.89 119.72 ;
      RECT 232.69 119.92 232.89 121.2 ;
      RECT 232.69 121.4 232.89 122.16 ;
      RECT 232.69 122.36 232.89 123.12 ;
      RECT 232.69 123.32 232.89 124.6 ;
      RECT 232.69 124.8 232.89 125.56 ;
      RECT 232.69 125.76 232.89 126.52 ;
      RECT 232.69 126.72 232.89 128 ;
      RECT 232.69 128.2 232.89 128.96 ;
      RECT 232.69 129.16 232.89 129.92 ;
      RECT 232.69 130.12 232.89 131.4 ;
      RECT 232.69 131.6 232.89 132.36 ;
      RECT 232.69 132.56 232.89 133.32 ;
      RECT 232.69 133.52 232.89 134.8 ;
      RECT 232.69 135 232.89 135.76 ;
      RECT 232.69 135.96 232.89 136.72 ;
      RECT 232.69 136.92 232.89 138.2 ;
      RECT 232.69 138.4 232.89 139.16 ;
      RECT 232.69 139.36 232.89 140.12 ;
      RECT 232.69 140.32 232.89 141.6 ;
      RECT 232.69 141.8 232.89 142.56 ;
      RECT 232.69 142.76 232.89 143.52 ;
      RECT 232.69 143.72 232.89 145 ;
      RECT 232.69 145.2 232.89 145.96 ;
      RECT 232.69 146.16 232.89 146.92 ;
      RECT 232.69 147.12 232.89 148.4 ;
      RECT 232.69 148.6 232.89 149.36 ;
      RECT 232.69 149.56 232.89 150.32 ;
      RECT 232.69 150.52 232.89 151.8 ;
      RECT 232.69 152 232.89 152.76 ;
      RECT 232.69 152.96 232.89 153.72 ;
      RECT 232.69 153.92 232.89 155.2 ;
      RECT 232.69 155.4 232.89 156.16 ;
      RECT 232.69 156.36 232.89 157.12 ;
      RECT 232.69 157.32 232.89 158.6 ;
      RECT 232.69 158.8 232.89 159.56 ;
      RECT 232.69 159.76 232.89 160.52 ;
      RECT 232.69 160.72 232.89 162 ;
      RECT 232.69 162.2 232.89 162.96 ;
      RECT 232.69 163.16 232.89 163.92 ;
      RECT 232.69 164.12 232.89 165.4 ;
      RECT 232.69 165.6 232.89 166.36 ;
      RECT 232.69 166.56 232.89 167.32 ;
      RECT 232.69 167.52 232.89 168.8 ;
      RECT 232.69 169 232.89 169.76 ;
      RECT 232.69 169.96 232.89 170.72 ;
      RECT 232.69 170.92 232.89 172.2 ;
      RECT 232.69 172.4 232.89 173.16 ;
      RECT 232.69 173.36 232.89 174.12 ;
      RECT 232.69 174.32 232.89 175.6 ;
      RECT 232.69 175.8 232.89 176.56 ;
      RECT 232.69 176.76 232.89 177.52 ;
      RECT 232.69 177.72 232.89 179 ;
      RECT 232.69 179.2 232.89 179.96 ;
      RECT 232.69 180.16 232.89 180.92 ;
      RECT 232.69 181.12 232.89 182.4 ;
      RECT 232.69 182.6 232.89 183.36 ;
      RECT 232.69 183.56 232.89 184.32 ;
      RECT 232.69 184.52 232.89 185.8 ;
      RECT 232.69 186 232.89 186.76 ;
      RECT 232.69 186.96 232.89 187.72 ;
      RECT 232.69 187.92 232.89 189.2 ;
      RECT 232.69 189.4 232.89 190.16 ;
      RECT 232.69 190.36 232.89 191.12 ;
      RECT 232.69 191.32 232.89 192.6 ;
      RECT 232.69 192.8 232.89 193.56 ;
      RECT 232.69 193.76 232.89 194.52 ;
      RECT 232.69 194.72 232.89 196 ;
      RECT 232.69 196.2 232.89 196.96 ;
      RECT 232.69 197.16 232.89 197.92 ;
      RECT 232.69 198.12 232.89 199.4 ;
      RECT 232.69 199.6 232.89 200.36 ;
      RECT 232.69 200.56 232.89 201.32 ;
      RECT 232.69 201.52 232.89 202.8 ;
      RECT 232.69 203 232.89 203.76 ;
      RECT 232.69 203.96 232.89 204.72 ;
      RECT 232.69 204.92 232.89 206.2 ;
      RECT 232.69 206.4 232.89 207.16 ;
      RECT 232.69 207.36 232.89 208.12 ;
      RECT 232.69 208.32 232.89 209.6 ;
      RECT 232.69 209.8 232.89 210.56 ;
      RECT 232.69 210.76 232.89 211.52 ;
      RECT 232.69 211.72 232.89 213 ;
      RECT 232.69 213.2 232.89 213.96 ;
      RECT 232.69 214.16 232.89 214.92 ;
      RECT 232.69 215.12 232.89 216.4 ;
      RECT 232.69 216.6 232.89 217.36 ;
      RECT 232.69 217.56 232.89 218.32 ;
      RECT 232.69 218.52 232.89 219.8 ;
      RECT 232.69 220 232.89 220.76 ;
      RECT 232.69 220.96 232.89 221.72 ;
      RECT 232.69 221.92 232.89 223.2 ;
      RECT 232.69 223.4 232.89 224.16 ;
      RECT 232.69 224.36 232.89 225.12 ;
      RECT 232.69 225.32 232.89 226.6 ;
      RECT 232.69 226.8 232.89 227.56 ;
      RECT 232.69 227.76 232.89 228.52 ;
      RECT 232.69 228.72 232.89 230 ;
      RECT 232.69 230.2 232.89 230.96 ;
      RECT 232.69 231.16 232.89 231.92 ;
      RECT 232.69 232.12 232.89 233.4 ;
      RECT 232.69 233.6 232.89 234.36 ;
      RECT 232.69 234.56 232.89 235.32 ;
      RECT 232.69 235.52 232.89 236.8 ;
      RECT 232.69 237 232.89 237.76 ;
      RECT 232.69 237.96 232.89 238.72 ;
      RECT 232.69 238.92 232.89 240.2 ;
      RECT 232.69 240.4 232.89 241.16 ;
      RECT 232.69 241.36 232.89 242.12 ;
      RECT 232.69 242.32 232.89 243.6 ;
      RECT 232.69 243.8 232.89 244.56 ;
      RECT 232.69 244.76 232.89 245.52 ;
      RECT 232.69 245.72 232.89 247 ;
      RECT 232.69 247.2 232.89 247.96 ;
      RECT 232.69 248.16 232.89 248.92 ;
      RECT 232.69 249.12 232.89 250.4 ;
      RECT 232.69 250.6 232.89 251.36 ;
      RECT 232.69 251.56 232.89 252.32 ;
      RECT 232.69 252.52 232.89 253.8 ;
      RECT 232.69 254 232.89 254.76 ;
      RECT 232.69 254.96 232.89 255.72 ;
      RECT 232.69 255.92 232.89 257.2 ;
      RECT 232.69 257.4 232.89 258.16 ;
      RECT 232.69 258.36 232.89 259.12 ;
      RECT 232.69 259.32 232.89 260.6 ;
      RECT 232.69 260.8 232.89 261.56 ;
      RECT 232.69 261.76 232.89 262.52 ;
      RECT 232.69 262.72 232.89 264 ;
      RECT 232.69 264.2 232.89 264.96 ;
      RECT 232.69 265.16 232.89 265.92 ;
      RECT 232.69 266.12 232.89 267.4 ;
      RECT 232.69 267.6 232.89 268.36 ;
      RECT 232.69 268.56 232.89 269.32 ;
      RECT 232.69 269.52 232.89 270.8 ;
      RECT 232.69 271 232.89 271.76 ;
      RECT 232.69 271.96 232.89 272.72 ;
      RECT 232.69 272.92 232.89 274.2 ;
      RECT 232.69 274.4 232.89 275.16 ;
      RECT 232.69 275.36 232.89 276.12 ;
      RECT 232.69 276.32 232.89 277.6 ;
      RECT 232.69 277.8 232.89 278.56 ;
      RECT 232.69 278.76 232.89 279.52 ;
      RECT 232.69 279.72 232.89 281 ;
      RECT 232.69 281.2 232.89 281.96 ;
      RECT 232.69 282.16 232.89 282.92 ;
      RECT 232.69 283.12 232.89 284.4 ;
      RECT 232.69 284.6 232.89 285.36 ;
      RECT 232.69 285.56 232.89 286.32 ;
      RECT 232.69 286.52 232.89 287.8 ;
      RECT 232.69 288 232.89 288.76 ;
      RECT 232.69 288.96 232.89 289.72 ;
      RECT 232.69 289.92 232.89 291.2 ;
      RECT 232.69 291.4 232.89 292.16 ;
      RECT 232.69 292.36 232.89 293.12 ;
      RECT 232.69 293.32 232.89 294.6 ;
      RECT 232.69 294.8 232.89 295.56 ;
      RECT 232.69 295.76 232.89 296.52 ;
      RECT 232.69 296.72 232.89 298 ;
      RECT 232.69 298.2 232.89 298.96 ;
      RECT 232.69 299.16 232.89 299.92 ;
      RECT 232.69 300.12 232.89 301.4 ;
      RECT 232.69 301.6 232.89 302.36 ;
      RECT 232.69 302.56 232.89 303.32 ;
      RECT 232.69 303.52 232.89 304.8 ;
      RECT 232.69 305 232.89 305.76 ;
      RECT 232.69 305.96 232.89 306.72 ;
      RECT 232.69 306.92 232.89 308.2 ;
      RECT 232.69 308.4 232.89 309.16 ;
      RECT 232.69 309.36 232.89 310.12 ;
      RECT 232.69 310.32 232.89 311.6 ;
      RECT 232.69 311.8 232.89 312.56 ;
      RECT 232.69 312.76 232.89 313.52 ;
      RECT 232.69 313.72 232.89 315 ;
      RECT 232.69 315.2 232.89 315.96 ;
      RECT 232.69 316.16 232.89 316.92 ;
      RECT 232.69 317.12 232.89 318.4 ;
      RECT 232.69 318.6 232.89 319.36 ;
      RECT 232.69 319.56 232.89 320.32 ;
      RECT 232.69 320.52 232.89 321.8 ;
      RECT 232.69 322 232.89 322.76 ;
      RECT 232.69 322.96 232.89 323.72 ;
      RECT 232.69 323.92 232.89 325.2 ;
      RECT 232.69 325.4 232.89 326.16 ;
      RECT 232.69 326.36 232.89 327.12 ;
      RECT 232.69 327.32 232.89 328.6 ;
      RECT 232.69 328.8 232.89 329.56 ;
      RECT 232.69 329.76 232.89 330.52 ;
      RECT 232.69 330.72 232.89 332 ;
      RECT 232.69 332.2 232.89 332.96 ;
      RECT 232.69 333.16 232.89 333.92 ;
      RECT 232.69 334.12 232.89 335.4 ;
      RECT 232.69 335.6 232.89 336.36 ;
      RECT 232.69 336.56 232.89 337.32 ;
      RECT 232.69 337.52 232.89 338.8 ;
      RECT 232.69 339 232.89 339.76 ;
      RECT 232.69 339.96 232.89 340.72 ;
      RECT 232.69 340.92 232.89 342.2 ;
      RECT 232.69 342.4 232.89 343.16 ;
      RECT 232.69 343.36 232.89 344.12 ;
      RECT 232.69 344.32 232.89 345.6 ;
      RECT 232.69 345.8 232.89 346.56 ;
      RECT 232.69 346.76 232.89 347.52 ;
      RECT 232.69 347.72 232.89 349 ;
      RECT 232.69 349.2 232.89 349.96 ;
      RECT 232.69 350.16 232.89 350.92 ;
      RECT 232.69 351.12 232.89 352.4 ;
      RECT 232.69 352.6 232.89 353.36 ;
      RECT 232.69 353.56 232.89 354.32 ;
      RECT 232.69 354.52 232.89 355.8 ;
      RECT 232.69 356 232.89 356.76 ;
      RECT 232.69 356.96 232.89 357.72 ;
      RECT 232.69 357.92 232.89 359.2 ;
      RECT 232.69 359.4 232.89 360.16 ;
      RECT 232.69 360.36 232.89 361.12 ;
      RECT 232.69 361.32 232.89 362.6 ;
      RECT 232.69 362.8 232.89 363.56 ;
      RECT 232.69 363.76 232.89 364.52 ;
      RECT 232.69 364.72 232.89 366 ;
      RECT 232.69 366.2 232.89 366.96 ;
      RECT 232.69 367.16 232.89 367.92 ;
      RECT 232.69 368.12 232.89 369.4 ;
      RECT 232.69 369.6 232.89 370.36 ;
      RECT 232.69 370.56 232.89 371.32 ;
      RECT 232.69 371.52 232.89 372.8 ;
      RECT 232.69 373 232.89 373.76 ;
      RECT 232.69 373.96 232.89 374.72 ;
      RECT 232.69 374.92 232.89 376.2 ;
      RECT 232.69 376.4 232.89 377.16 ;
      RECT 232.69 377.36 232.89 378.12 ;
      RECT 232.69 378.32 232.89 379.6 ;
      RECT 232.69 379.8 232.89 380.56 ;
      RECT 232.69 380.76 232.89 381.52 ;
      RECT 232.69 381.72 232.89 383 ;
      RECT 232.69 383.2 232.89 383.96 ;
      RECT 232.69 384.16 232.89 384.92 ;
      RECT 232.69 385.12 232.89 386.4 ;
      RECT 232.69 386.6 232.89 387.36 ;
      RECT 232.69 387.56 232.89 388.32 ;
      RECT 232.69 388.52 232.89 389.8 ;
      RECT 232.69 390 232.89 390.76 ;
      RECT 232.69 390.96 232.89 391.72 ;
      RECT 232.69 391.92 232.89 393.2 ;
      RECT 232.69 393.4 232.89 394.16 ;
      RECT 232.69 394.36 232.89 395.12 ;
      RECT 232.69 395.32 232.89 396.6 ;
      RECT 232.69 396.8 232.89 397.56 ;
      RECT 232.69 397.76 232.89 398.52 ;
      RECT 232.69 398.72 232.89 400 ;
      RECT 232.69 400.2 232.89 400.96 ;
      RECT 232.69 401.16 232.89 401.92 ;
      RECT 232.69 402.12 232.89 403.4 ;
      RECT 232.69 403.6 232.89 404.36 ;
      RECT 232.69 404.56 232.89 405.32 ;
      RECT 232.69 405.52 232.89 406.8 ;
      RECT 232.69 407 232.89 407.76 ;
      RECT 232.69 407.96 232.89 408.72 ;
      RECT 232.69 408.92 232.89 410.2 ;
      RECT 232.69 410.4 232.89 411.16 ;
      RECT 232.69 411.36 232.89 412.12 ;
      RECT 232.69 412.32 232.89 413.6 ;
      RECT 232.69 413.8 232.89 414.56 ;
      RECT 232.69 414.76 232.89 415.52 ;
      RECT 232.69 415.72 232.89 417 ;
      RECT 232.69 417.2 232.89 417.96 ;
      RECT 232.69 418.16 232.89 418.92 ;
      RECT 232.69 419.12 232.89 420.4 ;
      RECT 232.69 420.6 232.89 421.36 ;
      RECT 232.69 421.56 232.89 422.32 ;
      RECT 232.69 422.52 232.89 423.8 ;
      RECT 232.69 424 232.89 424.76 ;
      RECT 232.69 424.96 232.89 425.72 ;
      RECT 232.69 425.92 232.89 427.2 ;
      RECT 232.69 427.4 232.89 428.16 ;
      RECT 232.69 428.36 232.89 429.12 ;
      RECT 232.69 429.32 232.89 430.6 ;
      RECT 232.69 430.8 232.89 431.56 ;
      RECT 232.69 431.76 232.89 432.52 ;
      RECT 232.69 432.72 232.89 434 ;
      RECT 232.69 434.2 232.89 434.96 ;
      RECT 232.69 435.16 232.89 435.92 ;
      RECT 232.69 436.12 232.89 437.4 ;
      RECT 232.69 437.6 232.89 438.36 ;
      RECT 232.69 438.56 232.89 439.32 ;
      RECT 232.69 439.52 232.89 440.8 ;
      RECT 232.69 441 232.89 441.76 ;
      RECT 232.69 441.96 232.89 442.72 ;
      RECT 232.69 442.92 232.89 444.2 ;
      RECT 232.69 444.4 232.89 445.16 ;
      RECT 232.69 445.36 232.89 446.12 ;
      RECT 232.69 446.32 232.89 447.6 ;
      RECT 232.69 447.8 232.89 448.56 ;
      RECT 232.69 448.76 232.89 449.52 ;
      RECT 232.69 449.72 232.89 451 ;
      RECT 232.69 451.2 232.89 451.96 ;
      RECT 232.69 452.16 232.89 452.92 ;
      RECT 232.69 453.12 232.89 454.4 ;
      RECT 232.69 454.6 232.89 455.36 ;
      RECT 232.69 455.56 232.89 456.32 ;
      RECT 232.69 456.52 232.89 457.8 ;
      RECT 232.69 458 232.89 458.76 ;
      RECT 232.69 458.96 232.89 459.72 ;
      RECT 232.69 459.92 232.89 461.2 ;
      RECT 232.69 461.4 232.89 462.16 ;
      RECT 232.69 462.36 232.89 463.12 ;
      RECT 232.69 463.32 232.89 464.6 ;
      RECT 232.69 464.8 232.89 465.56 ;
      RECT 232.69 465.76 232.89 466.52 ;
      RECT 232.69 466.72 232.89 468 ;
      RECT 232.69 468.2 232.89 468.96 ;
      RECT 232.69 469.16 232.89 469.92 ;
      RECT 232.69 470.12 232.89 471.4 ;
      RECT 232.69 471.6 232.89 472.36 ;
      RECT 232.69 472.56 232.89 473.32 ;
      RECT 232.69 473.52 232.89 474.8 ;
      RECT 232.69 475 232.89 475.76 ;
      RECT 232.69 475.96 232.89 476.72 ;
      RECT 232.69 476.92 232.89 478.2 ;
      RECT 232.69 478.4 232.89 479.16 ;
      RECT 232.69 479.36 232.89 480.12 ;
      RECT 232.69 480.32 232.89 481.6 ;
      RECT 232.69 481.8 232.89 482.56 ;
      RECT 232.69 482.76 232.89 483.52 ;
      RECT 232.69 483.72 232.89 485 ;
      RECT 232.69 485.2 232.89 485.96 ;
      RECT 232.69 486.16 232.89 486.92 ;
      RECT 232.69 487.12 232.89 488.4 ;
      RECT 232.69 488.6 232.89 489.36 ;
      RECT 232.69 489.56 232.89 490.32 ;
      RECT 232.69 490.52 232.89 491.8 ;
      RECT 232.69 492 232.89 492.76 ;
      RECT 232.69 492.96 232.89 493.72 ;
      RECT 232.69 493.92 232.89 495.2 ;
      RECT 232.69 495.4 232.89 496.16 ;
      RECT 232.69 496.36 232.89 497.12 ;
      RECT 232.69 497.32 232.89 498.6 ;
      RECT 232.69 498.8 232.89 499.56 ;
      RECT 232.69 499.76 232.89 500.52 ;
      RECT 232.69 500.72 232.89 502 ;
      RECT 232.69 502.2 232.89 502.96 ;
      RECT 232.69 503.16 232.89 503.92 ;
      RECT 232.69 504.12 232.89 506.44 ;
      RECT 232.69 506.64 232.89 507.4 ;
      RECT 232.69 507.6 232.89 508.36 ;
      RECT 232.69 508.56 232.89 510 ;
      RECT 7.91 44.24 232.69 44.54 ;
      RECT 7.91 44.84 232.69 45.14 ;
      RECT 7.91 45.44 232.69 45.74 ;
      RECT 7.91 46.04 232.69 46.34 ;
      RECT 7.91 46.64 232.69 46.94 ;
      RECT 7.91 47.24 232.69 47.54 ;
      RECT 7.91 47.84 232.69 48.14 ;
      RECT 7.91 48.44 232.69 48.74 ;
      RECT 7.91 49.04 232.69 49.34 ;
      RECT 7.91 49.64 232.69 49.94 ;
      RECT 152.09 52.04 232.39 52.84 ;
      RECT 8.31 7.64 232.29 7.84 ;
      RECT 231.89 505.38 232.09 510.01 ;
      RECT 231.29 35.31 231.89 35.51 ;
      RECT 231.37 30.13 231.69 30.73 ;
      RECT 231.37 42.75 231.69 43.35 ;
      RECT 223.29 28.15 231.49 28.75 ;
      RECT 230.69 59.37 231.33 59.97 ;
      RECT 212.39 35.75 231.29 35.95 ;
      RECT 212.39 37.21 231.29 37.41 ;
      RECT 231.09 63.99 231.29 505.18 ;
      RECT 231.09 505.38 231.29 510.01 ;
      RECT 212.39 34.65 231.09 34.85 ;
      RECT 230.69 505.38 230.89 510.01 ;
      RECT 228.81 6.24 230.79 6.84 ;
      RECT 230.09 35.31 230.69 35.51 ;
      RECT 230.29 30.13 230.61 30.73 ;
      RECT 230.29 42.75 230.61 43.35 ;
      RECT 229.89 505.38 230.09 510.01 ;
      RECT 229.49 505.38 229.69 510.01 ;
      RECT 228.89 35.31 229.49 35.51 ;
      RECT 228.97 30.13 229.29 30.73 ;
      RECT 228.97 42.75 229.29 43.35 ;
      RECT 229.09 65.96 229.29 510.01 ;
      RECT 228.25 59.37 228.89 59.97 ;
      RECT 228.69 505.38 228.89 510.01 ;
      RECT 228.29 63.99 228.49 505.18 ;
      RECT 228.29 505.38 228.49 510.01 ;
      RECT 226.41 6.24 228.39 6.84 ;
      RECT 227.69 35.31 228.29 35.51 ;
      RECT 227.89 30.13 228.21 30.73 ;
      RECT 227.89 42.75 228.21 43.35 ;
      RECT 226.69 15.51 228.09 15.71 ;
      RECT 227.89 65.96 228.09 510.01 ;
      RECT 227.49 505.38 227.69 510.01 ;
      RECT 227.09 505.38 227.29 510.01 ;
      RECT 226.49 35.31 227.09 35.51 ;
      RECT 226.57 30.13 226.89 30.73 ;
      RECT 226.57 42.75 226.89 43.35 ;
      RECT 225.89 59.37 226.53 59.97 ;
      RECT 226.29 63.99 226.49 505.18 ;
      RECT 226.29 505.38 226.49 510.01 ;
      RECT 225.89 505.38 226.09 510.01 ;
      RECT 224.01 6.24 225.99 6.84 ;
      RECT 225.29 35.31 225.89 35.51 ;
      RECT 225.49 30.13 225.81 30.73 ;
      RECT 225.49 42.75 225.81 43.35 ;
      RECT 225.09 505.38 225.29 510.01 ;
      RECT 224.69 505.38 224.89 510.01 ;
      RECT 224.09 35.31 224.69 35.51 ;
      RECT 224.17 30.13 224.49 30.73 ;
      RECT 224.17 42.75 224.49 43.35 ;
      RECT 224.29 65.96 224.49 510.01 ;
      RECT 223.45 59.37 224.09 59.97 ;
      RECT 223.89 505.38 224.09 510.01 ;
      RECT 223.49 63.99 223.69 505.18 ;
      RECT 223.49 505.38 223.69 510.01 ;
      RECT 221.59 6.24 223.59 6.84 ;
      RECT 222.89 35.31 223.49 35.51 ;
      RECT 223.09 30.13 223.41 30.73 ;
      RECT 223.09 42.75 223.41 43.35 ;
      RECT 223.09 65.96 223.29 510.01 ;
      RECT 222.43 12.98 223.03 13.18 ;
      RECT 222.69 505.38 222.89 510.01 ;
      RECT 222.29 505.38 222.49 510.01 ;
      RECT 221.33 8.94 222.29 9.14 ;
      RECT 221.69 35.31 222.29 35.51 ;
      RECT 217.83 13.78 222.19 13.98 ;
      RECT 221.77 30.13 222.09 30.73 ;
      RECT 221.77 42.75 222.09 43.35 ;
      RECT 221.74 28.03 221.94 28.77 ;
      RECT 213.79 21.31 221.79 21.51 ;
      RECT 219.83 20.61 221.78 21.01 ;
      RECT 221.09 59.37 221.73 59.97 ;
      RECT 221.49 63.99 221.69 505.18 ;
      RECT 221.49 505.38 221.69 510.01 ;
      RECT 18.94 7.04 221.68 7.24 ;
      RECT 220.5 16.58 221.54 16.78 ;
      RECT 214.04 27.51 221.54 27.71 ;
      RECT 214.04 27.91 221.54 28.11 ;
      RECT 221.09 505.38 221.29 510.01 ;
      RECT 219.21 6.24 221.19 6.84 ;
      RECT 220.49 35.31 221.09 35.51 ;
      RECT 214.51 22.31 221.07 22.51 ;
      RECT 220.69 30.13 221.01 30.73 ;
      RECT 220.69 42.75 221.01 43.35 ;
      RECT 214.75 9.98 220.87 10.18 ;
      RECT 219.75 23.11 220.79 23.31 ;
      RECT 213.49 13.38 220.67 13.58 ;
      RECT 219.89 28.72 220.49 28.92 ;
      RECT 220.29 505.38 220.49 510.01 ;
      RECT 219.75 8.94 220.35 9.14 ;
      RECT 219.89 505.38 220.09 510.01 ;
      RECT 218.98 15.39 220.06 15.59 ;
      RECT 215.63 28.31 219.95 28.51 ;
      RECT 219.29 35.31 219.89 35.51 ;
      RECT 219.19 12.98 219.79 13.18 ;
      RECT 219.37 30.13 219.69 30.73 ;
      RECT 219.37 42.75 219.69 43.35 ;
      RECT 219.49 65.96 219.69 510.01 ;
      RECT 219.33 24.3 219.53 25.07 ;
      RECT 216.13 20.79 219.45 20.99 ;
      RECT 218.65 59.37 219.29 59.97 ;
      RECT 219.09 505.38 219.29 510.01 ;
      RECT 217.19 8.94 218.91 9.14 ;
      RECT 218.69 63.99 218.89 505.18 ;
      RECT 218.69 505.38 218.89 510.01 ;
      RECT 217.29 6.24 218.79 6.84 ;
      RECT 218.09 35.31 218.69 35.51 ;
      RECT 218.29 30.13 218.61 30.73 ;
      RECT 218.29 42.75 218.61 43.35 ;
      RECT 218.29 65.96 218.49 510.01 ;
      RECT 217.39 15.38 218.39 15.72 ;
      RECT 217.23 20.38 218.35 20.58 ;
      RECT 217.89 505.38 218.09 510.01 ;
      RECT 217.49 505.38 217.69 510.01 ;
      RECT 216.89 35.31 217.49 35.51 ;
      RECT 216.97 30.13 217.29 30.73 ;
      RECT 216.97 42.75 217.29 43.35 ;
      RECT 213.39 16.5 217.25 16.7 ;
      RECT 215.39 15.38 217.07 15.58 ;
      RECT 216.39 8.94 216.99 9.14 ;
      RECT 216.29 59.37 216.93 59.97 ;
      RECT 216.69 63.99 216.89 505.18 ;
      RECT 216.69 505.38 216.89 510.01 ;
      RECT 216.29 505.38 216.49 510.01 ;
      RECT 214.87 12.58 216.29 12.78 ;
      RECT 215.69 35.31 216.29 35.51 ;
      RECT 216.05 24.3 216.25 25.07 ;
      RECT 215.89 30.13 216.21 30.73 ;
      RECT 215.89 42.75 216.21 43.35 ;
      RECT 215.39 18.61 215.99 18.81 ;
      RECT 214.89 6.24 215.89 6.84 ;
      RECT 214.79 23.11 215.83 23.31 ;
      RECT 213.8 20.61 215.75 21.01 ;
      RECT 215.09 28.72 215.69 28.92 ;
      RECT 215.49 505.38 215.69 510.01 ;
      RECT 215.09 505.38 215.29 510.01 ;
      RECT 214.49 35.31 215.09 35.51 ;
      RECT 214.57 30.13 214.89 30.73 ;
      RECT 214.57 42.75 214.89 43.35 ;
      RECT 214.69 65.96 214.89 510.01 ;
      RECT 213.85 59.37 214.49 59.97 ;
      RECT 214.29 505.38 214.49 510.01 ;
      RECT 213.89 63.99 214.09 505.18 ;
      RECT 213.89 505.38 214.09 510.01 ;
      RECT 213.29 35.31 213.89 35.51 ;
      RECT 213.64 28.03 213.84 28.77 ;
      RECT 213.49 30.13 213.81 30.73 ;
      RECT 213.49 42.75 213.81 43.35 ;
      RECT 213.49 65.96 213.69 510.01 ;
      RECT 213.39 15.38 213.59 15.98 ;
      RECT 212.59 6.24 213.39 6.84 ;
      RECT 213.09 505.38 213.29 510.01 ;
      RECT 212.89 12.58 213.09 13.85 ;
      RECT 212.69 505.38 212.89 510.01 ;
      RECT 212.09 35.31 212.69 35.51 ;
      RECT 212.39 15.38 212.59 15.98 ;
      RECT 208.73 16.5 212.59 16.7 ;
      RECT 205.31 13.38 212.49 13.58 ;
      RECT 212.17 30.13 212.49 30.73 ;
      RECT 212.17 42.75 212.49 43.35 ;
      RECT 212.14 28.03 212.34 28.77 ;
      RECT 204.19 21.31 212.19 21.51 ;
      RECT 210.23 20.61 212.18 21.01 ;
      RECT 211.49 59.37 212.13 59.97 ;
      RECT 191.99 35.75 212.09 35.95 ;
      RECT 191.99 37.21 212.09 37.41 ;
      RECT 211.89 63.99 212.09 505.18 ;
      RECT 211.89 505.38 212.09 510.01 ;
      RECT 204.44 27.51 211.94 27.71 ;
      RECT 204.44 27.91 211.94 28.11 ;
      RECT 191.99 34.65 211.89 34.85 ;
      RECT 211.49 505.38 211.69 510.01 ;
      RECT 210.89 35.31 211.49 35.51 ;
      RECT 204.91 22.31 211.47 22.51 ;
      RECT 211.09 30.13 211.41 30.73 ;
      RECT 211.09 42.75 211.41 43.35 ;
      RECT 205.11 9.98 211.23 10.18 ;
      RECT 210.15 23.11 211.19 23.31 ;
      RECT 209.69 12.58 211.11 12.78 ;
      RECT 210.09 6.24 211.09 6.84 ;
      RECT 210.29 28.72 210.89 28.92 ;
      RECT 210.69 505.38 210.89 510.01 ;
      RECT 208.91 15.38 210.59 15.58 ;
      RECT 209.99 18.61 210.59 18.81 ;
      RECT 210.29 505.38 210.49 510.01 ;
      RECT 206.03 28.31 210.35 28.51 ;
      RECT 209.69 35.31 210.29 35.51 ;
      RECT 209.77 30.13 210.09 30.73 ;
      RECT 209.77 42.75 210.09 43.35 ;
      RECT 209.89 65.96 210.09 510.01 ;
      RECT 209.73 24.3 209.93 25.07 ;
      RECT 206.53 20.79 209.85 20.99 ;
      RECT 209.05 59.37 209.69 59.97 ;
      RECT 209.49 505.38 209.69 510.01 ;
      RECT 208.99 8.94 209.59 9.14 ;
      RECT 209.09 63.99 209.29 505.18 ;
      RECT 209.09 505.38 209.29 510.01 ;
      RECT 208.49 35.31 209.09 35.51 ;
      RECT 208.69 30.13 209.01 30.73 ;
      RECT 208.69 42.75 209.01 43.35 ;
      RECT 208.69 65.96 208.89 510.01 ;
      RECT 207.07 8.94 208.79 9.14 ;
      RECT 207.63 20.38 208.75 20.58 ;
      RECT 207.19 6.24 208.69 6.84 ;
      RECT 207.59 15.38 208.59 15.72 ;
      RECT 208.29 505.38 208.49 510.01 ;
      RECT 203.79 13.78 208.15 13.98 ;
      RECT 207.89 505.38 208.09 510.01 ;
      RECT 207.29 35.31 207.89 35.51 ;
      RECT 207.37 30.13 207.69 30.73 ;
      RECT 207.37 42.75 207.69 43.35 ;
      RECT 206.69 59.37 207.33 59.97 ;
      RECT 207.09 63.99 207.29 505.18 ;
      RECT 207.09 505.38 207.29 510.01 ;
      RECT 205.92 15.39 207 15.59 ;
      RECT 206.69 505.38 206.89 510.01 ;
      RECT 206.19 12.98 206.79 13.18 ;
      RECT 204.79 6.24 206.76 6.84 ;
      RECT 206.09 35.31 206.69 35.51 ;
      RECT 206.45 24.3 206.65 25.07 ;
      RECT 206.29 30.13 206.61 30.73 ;
      RECT 206.29 42.75 206.61 43.35 ;
      RECT 205.63 8.94 206.23 9.14 ;
      RECT 205.19 23.11 206.23 23.31 ;
      RECT 204.2 20.61 206.15 21.01 ;
      RECT 205.49 28.72 206.09 28.92 ;
      RECT 205.89 505.38 206.09 510.01 ;
      RECT 205.49 505.38 205.69 510.01 ;
      RECT 204.89 35.31 205.49 35.51 ;
      RECT 204.44 16.58 205.48 16.78 ;
      RECT 204.97 30.13 205.29 30.73 ;
      RECT 204.97 42.75 205.29 43.35 ;
      RECT 205.09 65.96 205.29 510.01 ;
      RECT 204.25 59.37 204.89 59.97 ;
      RECT 204.69 505.38 204.89 510.01 ;
      RECT 203.69 8.94 204.65 9.14 ;
      RECT 204.29 63.99 204.49 505.18 ;
      RECT 204.29 505.38 204.49 510.01 ;
      RECT 202.39 6.24 204.39 6.84 ;
      RECT 203.69 35.31 204.29 35.51 ;
      RECT 204.04 28.03 204.24 28.77 ;
      RECT 203.89 30.13 204.21 30.73 ;
      RECT 203.89 42.75 204.21 43.35 ;
      RECT 203.89 65.96 204.09 510.01 ;
      RECT 203.49 505.38 203.69 510.01 ;
      RECT 202.95 12.98 203.55 13.18 ;
      RECT 203.09 505.38 203.29 510.01 ;
      RECT 202.49 35.31 203.09 35.51 ;
      RECT 202.57 30.13 202.89 30.73 ;
      RECT 202.57 42.75 202.89 43.35 ;
      RECT 194.49 28.15 202.69 28.75 ;
      RECT 201.89 59.37 202.53 59.97 ;
      RECT 202.29 63.99 202.49 505.18 ;
      RECT 202.29 505.38 202.49 510.01 ;
      RECT 201.89 505.38 202.09 510.01 ;
      RECT 199.99 6.24 201.97 6.84 ;
      RECT 201.29 35.31 201.89 35.51 ;
      RECT 201.49 30.13 201.81 30.73 ;
      RECT 201.49 42.75 201.81 43.35 ;
      RECT 201.09 505.38 201.29 510.01 ;
      RECT 200.69 505.38 200.89 510.01 ;
      RECT 200.09 35.31 200.69 35.51 ;
      RECT 200.17 30.13 200.49 30.73 ;
      RECT 200.17 42.75 200.49 43.35 ;
      RECT 200.29 65.96 200.49 510.01 ;
      RECT 199.45 59.37 200.09 59.97 ;
      RECT 199.89 505.38 200.09 510.01 ;
      RECT 199.49 63.99 199.69 505.18 ;
      RECT 199.49 505.38 199.69 510.01 ;
      RECT 197.59 6.24 199.57 6.84 ;
      RECT 198.89 35.31 199.49 35.51 ;
      RECT 199.09 30.13 199.41 30.73 ;
      RECT 199.09 42.75 199.41 43.35 ;
      RECT 197.89 15.51 199.29 15.71 ;
      RECT 199.09 65.96 199.29 510.01 ;
      RECT 198.69 505.38 198.89 510.01 ;
      RECT 198.29 505.38 198.49 510.01 ;
      RECT 197.69 35.31 198.29 35.51 ;
      RECT 197.77 30.13 198.09 30.73 ;
      RECT 197.77 42.75 198.09 43.35 ;
      RECT 197.09 59.37 197.73 59.97 ;
      RECT 197.49 63.99 197.69 505.18 ;
      RECT 197.49 505.38 197.69 510.01 ;
      RECT 197.09 505.38 197.29 510.01 ;
      RECT 195.19 6.24 197.17 6.84 ;
      RECT 196.49 35.31 197.09 35.51 ;
      RECT 196.69 30.13 197.01 30.73 ;
      RECT 196.69 42.75 197.01 43.35 ;
      RECT 196.29 505.38 196.49 510.01 ;
      RECT 195.89 505.38 196.09 510.01 ;
      RECT 195.29 35.31 195.89 35.51 ;
      RECT 195.37 30.13 195.69 30.73 ;
      RECT 195.37 42.75 195.69 43.35 ;
      RECT 195.49 65.96 195.69 510.01 ;
      RECT 194.65 59.37 195.29 59.97 ;
      RECT 195.09 505.38 195.29 510.01 ;
      RECT 194.69 63.99 194.89 505.18 ;
      RECT 194.69 505.38 194.89 510.01 ;
      RECT 193.39 6.24 194.79 6.84 ;
      RECT 194.09 35.31 194.69 35.51 ;
      RECT 194.29 30.13 194.61 30.73 ;
      RECT 194.29 42.75 194.61 43.35 ;
      RECT 194.29 65.96 194.49 510.01 ;
      RECT 193.89 505.38 194.09 510.01 ;
      RECT 193.09 68.76 193.29 70.14 ;
      RECT 193.09 70.34 193.29 71.16 ;
      RECT 193.09 71.36 193.29 72.18 ;
      RECT 193.09 72.38 193.29 73.54 ;
      RECT 193.09 73.74 193.29 74.56 ;
      RECT 193.09 74.76 193.29 75.58 ;
      RECT 193.09 75.78 193.29 76.94 ;
      RECT 193.09 77.14 193.29 77.96 ;
      RECT 193.09 78.16 193.29 78.98 ;
      RECT 193.09 79.18 193.29 80.34 ;
      RECT 193.09 80.54 193.29 81.36 ;
      RECT 193.09 81.56 193.29 82.38 ;
      RECT 193.09 82.58 193.29 83.74 ;
      RECT 193.09 83.94 193.29 84.76 ;
      RECT 193.09 84.96 193.29 85.78 ;
      RECT 193.09 85.98 193.29 87.14 ;
      RECT 193.09 87.34 193.29 88.16 ;
      RECT 193.09 88.36 193.29 89.18 ;
      RECT 193.09 89.38 193.29 90.54 ;
      RECT 193.09 90.74 193.29 91.56 ;
      RECT 193.09 91.76 193.29 92.58 ;
      RECT 193.09 92.78 193.29 93.94 ;
      RECT 193.09 94.14 193.29 94.96 ;
      RECT 193.09 95.16 193.29 95.98 ;
      RECT 193.09 96.18 193.29 97.34 ;
      RECT 193.09 97.54 193.29 98.36 ;
      RECT 193.09 98.56 193.29 99.38 ;
      RECT 193.09 99.58 193.29 100.74 ;
      RECT 193.09 100.94 193.29 101.76 ;
      RECT 193.09 101.96 193.29 102.78 ;
      RECT 193.09 102.98 193.29 104.14 ;
      RECT 193.09 104.34 193.29 105.16 ;
      RECT 193.09 105.36 193.29 106.18 ;
      RECT 193.09 106.38 193.29 107.54 ;
      RECT 193.09 107.74 193.29 108.56 ;
      RECT 193.09 108.76 193.29 109.58 ;
      RECT 193.09 109.78 193.29 110.94 ;
      RECT 193.09 111.14 193.29 111.96 ;
      RECT 193.09 112.16 193.29 112.98 ;
      RECT 193.09 113.18 193.29 114.34 ;
      RECT 193.09 114.54 193.29 115.36 ;
      RECT 193.09 115.56 193.29 116.38 ;
      RECT 193.09 116.58 193.29 117.74 ;
      RECT 193.09 117.94 193.29 118.76 ;
      RECT 193.09 118.96 193.29 119.78 ;
      RECT 193.09 119.98 193.29 121.14 ;
      RECT 193.09 121.34 193.29 122.16 ;
      RECT 193.09 122.36 193.29 123.18 ;
      RECT 193.09 123.38 193.29 124.54 ;
      RECT 193.09 124.74 193.29 125.56 ;
      RECT 193.09 125.76 193.29 126.58 ;
      RECT 193.09 126.78 193.29 127.94 ;
      RECT 193.09 128.14 193.29 128.96 ;
      RECT 193.09 129.16 193.29 129.98 ;
      RECT 193.09 130.18 193.29 131.34 ;
      RECT 193.09 131.54 193.29 132.36 ;
      RECT 193.09 132.56 193.29 133.38 ;
      RECT 193.09 133.58 193.29 134.74 ;
      RECT 193.09 134.94 193.29 135.76 ;
      RECT 193.09 135.96 193.29 136.78 ;
      RECT 193.09 136.98 193.29 138.14 ;
      RECT 193.09 138.34 193.29 139.16 ;
      RECT 193.09 139.36 193.29 140.18 ;
      RECT 193.09 140.38 193.29 141.54 ;
      RECT 193.09 141.74 193.29 142.56 ;
      RECT 193.09 142.76 193.29 143.58 ;
      RECT 193.09 143.78 193.29 144.94 ;
      RECT 193.09 145.14 193.29 145.96 ;
      RECT 193.09 146.16 193.29 146.98 ;
      RECT 193.09 147.18 193.29 148.34 ;
      RECT 193.09 148.54 193.29 149.36 ;
      RECT 193.09 149.56 193.29 150.38 ;
      RECT 193.09 150.58 193.29 151.74 ;
      RECT 193.09 151.94 193.29 152.76 ;
      RECT 193.09 152.96 193.29 153.78 ;
      RECT 193.09 153.98 193.29 155.14 ;
      RECT 193.09 155.34 193.29 156.16 ;
      RECT 193.09 156.36 193.29 157.18 ;
      RECT 193.09 157.38 193.29 158.54 ;
      RECT 193.09 158.74 193.29 159.56 ;
      RECT 193.09 159.76 193.29 160.58 ;
      RECT 193.09 160.78 193.29 161.94 ;
      RECT 193.09 162.14 193.29 162.96 ;
      RECT 193.09 163.16 193.29 163.98 ;
      RECT 193.09 164.18 193.29 165.34 ;
      RECT 193.09 165.54 193.29 166.36 ;
      RECT 193.09 166.56 193.29 167.38 ;
      RECT 193.09 167.58 193.29 168.74 ;
      RECT 193.09 168.94 193.29 169.76 ;
      RECT 193.09 169.96 193.29 170.78 ;
      RECT 193.09 170.98 193.29 172.14 ;
      RECT 193.09 172.34 193.29 173.16 ;
      RECT 193.09 173.36 193.29 174.18 ;
      RECT 193.09 174.38 193.29 175.54 ;
      RECT 193.09 175.74 193.29 176.56 ;
      RECT 193.09 176.76 193.29 177.58 ;
      RECT 193.09 177.78 193.29 178.94 ;
      RECT 193.09 179.14 193.29 179.96 ;
      RECT 193.09 180.16 193.29 180.98 ;
      RECT 193.09 181.18 193.29 182.34 ;
      RECT 193.09 182.54 193.29 183.36 ;
      RECT 193.09 183.56 193.29 184.38 ;
      RECT 193.09 184.58 193.29 185.74 ;
      RECT 193.09 185.94 193.29 186.76 ;
      RECT 193.09 186.96 193.29 187.78 ;
      RECT 193.09 187.98 193.29 189.14 ;
      RECT 193.09 189.34 193.29 190.16 ;
      RECT 193.09 190.36 193.29 191.18 ;
      RECT 193.09 191.38 193.29 192.54 ;
      RECT 193.09 192.74 193.29 193.56 ;
      RECT 193.09 193.76 193.29 194.58 ;
      RECT 193.09 194.78 193.29 195.94 ;
      RECT 193.09 196.14 193.29 196.96 ;
      RECT 193.09 197.16 193.29 197.98 ;
      RECT 193.09 198.18 193.29 199.34 ;
      RECT 193.09 199.54 193.29 200.36 ;
      RECT 193.09 200.56 193.29 201.38 ;
      RECT 193.09 201.58 193.29 202.74 ;
      RECT 193.09 202.94 193.29 203.76 ;
      RECT 193.09 203.96 193.29 204.78 ;
      RECT 193.09 204.98 193.29 206.14 ;
      RECT 193.09 206.34 193.29 207.16 ;
      RECT 193.09 207.36 193.29 208.18 ;
      RECT 193.09 208.38 193.29 209.54 ;
      RECT 193.09 209.74 193.29 210.56 ;
      RECT 193.09 210.76 193.29 211.58 ;
      RECT 193.09 211.78 193.29 212.94 ;
      RECT 193.09 213.14 193.29 213.96 ;
      RECT 193.09 214.16 193.29 214.98 ;
      RECT 193.09 215.18 193.29 216.34 ;
      RECT 193.09 216.54 193.29 217.36 ;
      RECT 193.09 217.56 193.29 218.38 ;
      RECT 193.09 218.58 193.29 219.74 ;
      RECT 193.09 219.94 193.29 220.76 ;
      RECT 193.09 220.96 193.29 221.78 ;
      RECT 193.09 221.98 193.29 223.14 ;
      RECT 193.09 223.34 193.29 224.16 ;
      RECT 193.09 224.36 193.29 225.18 ;
      RECT 193.09 225.38 193.29 226.54 ;
      RECT 193.09 226.74 193.29 227.56 ;
      RECT 193.09 227.76 193.29 228.58 ;
      RECT 193.09 228.78 193.29 229.94 ;
      RECT 193.09 230.14 193.29 230.96 ;
      RECT 193.09 231.16 193.29 231.98 ;
      RECT 193.09 232.18 193.29 233.34 ;
      RECT 193.09 233.54 193.29 234.36 ;
      RECT 193.09 234.56 193.29 235.38 ;
      RECT 193.09 235.58 193.29 236.74 ;
      RECT 193.09 236.94 193.29 237.76 ;
      RECT 193.09 237.96 193.29 238.78 ;
      RECT 193.09 238.98 193.29 240.14 ;
      RECT 193.09 240.34 193.29 241.16 ;
      RECT 193.09 241.36 193.29 242.18 ;
      RECT 193.09 242.38 193.29 243.54 ;
      RECT 193.09 243.74 193.29 244.56 ;
      RECT 193.09 244.76 193.29 245.58 ;
      RECT 193.09 245.78 193.29 246.94 ;
      RECT 193.09 247.14 193.29 247.96 ;
      RECT 193.09 248.16 193.29 248.98 ;
      RECT 193.09 249.18 193.29 250.34 ;
      RECT 193.09 250.54 193.29 251.36 ;
      RECT 193.09 251.56 193.29 252.38 ;
      RECT 193.09 252.58 193.29 253.74 ;
      RECT 193.09 253.94 193.29 254.76 ;
      RECT 193.09 254.96 193.29 255.78 ;
      RECT 193.09 255.98 193.29 257.14 ;
      RECT 193.09 257.34 193.29 258.16 ;
      RECT 193.09 258.36 193.29 259.18 ;
      RECT 193.09 259.38 193.29 260.54 ;
      RECT 193.09 260.74 193.29 261.56 ;
      RECT 193.09 261.76 193.29 262.58 ;
      RECT 193.09 262.78 193.29 263.94 ;
      RECT 193.09 264.14 193.29 264.96 ;
      RECT 193.09 265.16 193.29 265.98 ;
      RECT 193.09 266.18 193.29 267.34 ;
      RECT 193.09 267.54 193.29 268.36 ;
      RECT 193.09 268.56 193.29 269.38 ;
      RECT 193.09 269.58 193.29 270.74 ;
      RECT 193.09 270.94 193.29 271.76 ;
      RECT 193.09 271.96 193.29 272.78 ;
      RECT 193.09 272.98 193.29 274.14 ;
      RECT 193.09 274.34 193.29 275.16 ;
      RECT 193.09 275.36 193.29 276.18 ;
      RECT 193.09 276.38 193.29 277.54 ;
      RECT 193.09 277.74 193.29 278.56 ;
      RECT 193.09 278.76 193.29 279.58 ;
      RECT 193.09 279.78 193.29 280.94 ;
      RECT 193.09 281.14 193.29 281.96 ;
      RECT 193.09 282.16 193.29 282.98 ;
      RECT 193.09 283.18 193.29 284.34 ;
      RECT 193.09 284.54 193.29 285.36 ;
      RECT 193.09 285.56 193.29 286.38 ;
      RECT 193.09 286.58 193.29 287.74 ;
      RECT 193.09 287.94 193.29 288.76 ;
      RECT 193.09 288.96 193.29 289.78 ;
      RECT 193.09 289.98 193.29 291.14 ;
      RECT 193.09 291.34 193.29 292.16 ;
      RECT 193.09 292.36 193.29 293.18 ;
      RECT 193.09 293.38 193.29 294.54 ;
      RECT 193.09 294.74 193.29 295.56 ;
      RECT 193.09 295.76 193.29 296.58 ;
      RECT 193.09 296.78 193.29 297.94 ;
      RECT 193.09 298.14 193.29 298.96 ;
      RECT 193.09 299.16 193.29 299.98 ;
      RECT 193.09 300.18 193.29 301.34 ;
      RECT 193.09 301.54 193.29 302.36 ;
      RECT 193.09 302.56 193.29 303.38 ;
      RECT 193.09 303.58 193.29 304.74 ;
      RECT 193.09 304.94 193.29 305.76 ;
      RECT 193.09 305.96 193.29 306.78 ;
      RECT 193.09 306.98 193.29 308.14 ;
      RECT 193.09 308.34 193.29 309.16 ;
      RECT 193.09 309.36 193.29 310.18 ;
      RECT 193.09 310.38 193.29 311.54 ;
      RECT 193.09 311.74 193.29 312.56 ;
      RECT 193.09 312.76 193.29 313.58 ;
      RECT 193.09 313.78 193.29 314.94 ;
      RECT 193.09 315.14 193.29 315.96 ;
      RECT 193.09 316.16 193.29 316.98 ;
      RECT 193.09 317.18 193.29 318.34 ;
      RECT 193.09 318.54 193.29 319.36 ;
      RECT 193.09 319.56 193.29 320.38 ;
      RECT 193.09 320.58 193.29 321.74 ;
      RECT 193.09 321.94 193.29 322.76 ;
      RECT 193.09 322.96 193.29 323.78 ;
      RECT 193.09 323.98 193.29 325.14 ;
      RECT 193.09 325.34 193.29 326.16 ;
      RECT 193.09 326.36 193.29 327.18 ;
      RECT 193.09 327.38 193.29 328.54 ;
      RECT 193.09 328.74 193.29 329.56 ;
      RECT 193.09 329.76 193.29 330.58 ;
      RECT 193.09 330.78 193.29 331.94 ;
      RECT 193.09 332.14 193.29 332.96 ;
      RECT 193.09 333.16 193.29 333.98 ;
      RECT 193.09 334.18 193.29 335.34 ;
      RECT 193.09 335.54 193.29 336.36 ;
      RECT 193.09 336.56 193.29 337.38 ;
      RECT 193.09 337.58 193.29 338.74 ;
      RECT 193.09 338.94 193.29 339.76 ;
      RECT 193.09 339.96 193.29 340.78 ;
      RECT 193.09 340.98 193.29 342.14 ;
      RECT 193.09 342.34 193.29 343.16 ;
      RECT 193.09 343.36 193.29 344.18 ;
      RECT 193.09 344.38 193.29 345.54 ;
      RECT 193.09 345.74 193.29 346.56 ;
      RECT 193.09 346.76 193.29 347.58 ;
      RECT 193.09 347.78 193.29 348.94 ;
      RECT 193.09 349.14 193.29 349.96 ;
      RECT 193.09 350.16 193.29 350.98 ;
      RECT 193.09 351.18 193.29 352.34 ;
      RECT 193.09 352.54 193.29 353.36 ;
      RECT 193.09 353.56 193.29 354.38 ;
      RECT 193.09 354.58 193.29 355.74 ;
      RECT 193.09 355.94 193.29 356.76 ;
      RECT 193.09 356.96 193.29 357.78 ;
      RECT 193.09 357.98 193.29 359.14 ;
      RECT 193.09 359.34 193.29 360.16 ;
      RECT 193.09 360.36 193.29 361.18 ;
      RECT 193.09 361.38 193.29 362.54 ;
      RECT 193.09 362.74 193.29 363.56 ;
      RECT 193.09 363.76 193.29 364.58 ;
      RECT 193.09 364.78 193.29 365.94 ;
      RECT 193.09 366.14 193.29 366.96 ;
      RECT 193.09 367.16 193.29 367.98 ;
      RECT 193.09 368.18 193.29 369.34 ;
      RECT 193.09 369.54 193.29 370.36 ;
      RECT 193.09 370.56 193.29 371.38 ;
      RECT 193.09 371.58 193.29 372.74 ;
      RECT 193.09 372.94 193.29 373.76 ;
      RECT 193.09 373.96 193.29 374.78 ;
      RECT 193.09 374.98 193.29 376.14 ;
      RECT 193.09 376.34 193.29 377.16 ;
      RECT 193.09 377.36 193.29 378.18 ;
      RECT 193.09 378.38 193.29 379.54 ;
      RECT 193.09 379.74 193.29 380.56 ;
      RECT 193.09 380.76 193.29 381.58 ;
      RECT 193.09 381.78 193.29 382.94 ;
      RECT 193.09 383.14 193.29 383.96 ;
      RECT 193.09 384.16 193.29 384.98 ;
      RECT 193.09 385.18 193.29 386.34 ;
      RECT 193.09 386.54 193.29 387.36 ;
      RECT 193.09 387.56 193.29 388.38 ;
      RECT 193.09 388.58 193.29 389.74 ;
      RECT 193.09 389.94 193.29 390.76 ;
      RECT 193.09 390.96 193.29 391.78 ;
      RECT 193.09 391.98 193.29 393.14 ;
      RECT 193.09 393.34 193.29 394.16 ;
      RECT 193.09 394.36 193.29 395.18 ;
      RECT 193.09 395.38 193.29 396.54 ;
      RECT 193.09 396.74 193.29 397.56 ;
      RECT 193.09 397.76 193.29 398.58 ;
      RECT 193.09 398.78 193.29 399.94 ;
      RECT 193.09 400.14 193.29 400.96 ;
      RECT 193.09 401.16 193.29 401.98 ;
      RECT 193.09 402.18 193.29 403.34 ;
      RECT 193.09 403.54 193.29 404.36 ;
      RECT 193.09 404.56 193.29 405.38 ;
      RECT 193.09 405.58 193.29 406.74 ;
      RECT 193.09 406.94 193.29 407.76 ;
      RECT 193.09 407.96 193.29 408.78 ;
      RECT 193.09 408.98 193.29 410.14 ;
      RECT 193.09 410.34 193.29 411.16 ;
      RECT 193.09 411.36 193.29 412.18 ;
      RECT 193.09 412.38 193.29 413.54 ;
      RECT 193.09 413.74 193.29 414.56 ;
      RECT 193.09 414.76 193.29 415.58 ;
      RECT 193.09 415.78 193.29 416.94 ;
      RECT 193.09 417.14 193.29 417.96 ;
      RECT 193.09 418.16 193.29 418.98 ;
      RECT 193.09 419.18 193.29 420.34 ;
      RECT 193.09 420.54 193.29 421.36 ;
      RECT 193.09 421.56 193.29 422.38 ;
      RECT 193.09 422.58 193.29 423.74 ;
      RECT 193.09 423.94 193.29 424.76 ;
      RECT 193.09 424.96 193.29 425.78 ;
      RECT 193.09 425.98 193.29 427.14 ;
      RECT 193.09 427.34 193.29 428.16 ;
      RECT 193.09 428.36 193.29 429.18 ;
      RECT 193.09 429.38 193.29 430.54 ;
      RECT 193.09 430.74 193.29 431.56 ;
      RECT 193.09 431.76 193.29 432.58 ;
      RECT 193.09 432.78 193.29 433.94 ;
      RECT 193.09 434.14 193.29 434.96 ;
      RECT 193.09 435.16 193.29 435.98 ;
      RECT 193.09 436.18 193.29 437.34 ;
      RECT 193.09 437.54 193.29 438.36 ;
      RECT 193.09 438.56 193.29 439.38 ;
      RECT 193.09 439.58 193.29 440.74 ;
      RECT 193.09 440.94 193.29 441.76 ;
      RECT 193.09 441.96 193.29 442.78 ;
      RECT 193.09 442.98 193.29 444.14 ;
      RECT 193.09 444.34 193.29 445.16 ;
      RECT 193.09 445.36 193.29 446.18 ;
      RECT 193.09 446.38 193.29 447.54 ;
      RECT 193.09 447.74 193.29 448.56 ;
      RECT 193.09 448.76 193.29 449.58 ;
      RECT 193.09 449.78 193.29 450.94 ;
      RECT 193.09 451.14 193.29 451.96 ;
      RECT 193.09 452.16 193.29 452.98 ;
      RECT 193.09 453.18 193.29 454.34 ;
      RECT 193.09 454.54 193.29 455.36 ;
      RECT 193.09 455.56 193.29 456.38 ;
      RECT 193.09 456.58 193.29 457.74 ;
      RECT 193.09 457.94 193.29 458.76 ;
      RECT 193.09 458.96 193.29 459.78 ;
      RECT 193.09 459.98 193.29 461.14 ;
      RECT 193.09 461.34 193.29 462.16 ;
      RECT 193.09 462.36 193.29 463.18 ;
      RECT 193.09 463.38 193.29 464.54 ;
      RECT 193.09 464.74 193.29 465.56 ;
      RECT 193.09 465.76 193.29 466.58 ;
      RECT 193.09 466.78 193.29 467.94 ;
      RECT 193.09 468.14 193.29 468.96 ;
      RECT 193.09 469.16 193.29 469.98 ;
      RECT 193.09 470.18 193.29 471.34 ;
      RECT 193.09 471.54 193.29 472.36 ;
      RECT 193.09 472.56 193.29 473.38 ;
      RECT 193.09 473.58 193.29 474.74 ;
      RECT 193.09 474.94 193.29 475.76 ;
      RECT 193.09 475.96 193.29 476.78 ;
      RECT 193.09 476.98 193.29 478.14 ;
      RECT 193.09 478.34 193.29 479.16 ;
      RECT 193.09 479.36 193.29 480.18 ;
      RECT 193.09 480.38 193.29 481.54 ;
      RECT 193.09 481.74 193.29 482.56 ;
      RECT 193.09 482.76 193.29 483.58 ;
      RECT 193.09 483.78 193.29 484.94 ;
      RECT 193.09 485.14 193.29 485.96 ;
      RECT 193.09 486.16 193.29 486.98 ;
      RECT 193.09 487.18 193.29 488.34 ;
      RECT 193.09 488.54 193.29 489.36 ;
      RECT 193.09 489.56 193.29 490.38 ;
      RECT 193.09 490.58 193.29 491.74 ;
      RECT 193.09 491.94 193.29 492.76 ;
      RECT 193.09 492.96 193.29 493.78 ;
      RECT 193.09 493.98 193.29 495.14 ;
      RECT 193.09 495.34 193.29 496.16 ;
      RECT 193.09 496.36 193.29 497.18 ;
      RECT 193.09 497.38 193.29 498.54 ;
      RECT 193.09 498.74 193.29 499.56 ;
      RECT 193.09 499.76 193.29 500.58 ;
      RECT 193.09 500.78 193.29 501.94 ;
      RECT 193.09 502.14 193.29 502.96 ;
      RECT 193.09 503.16 193.29 503.98 ;
      RECT 193.09 504.18 193.29 506.38 ;
      RECT 193.09 506.58 193.29 507.4 ;
      RECT 193.09 507.6 193.29 508.42 ;
      RECT 193.09 508.62 193.29 510 ;
      RECT 191.59 6.24 192.99 6.84 ;
      RECT 192.29 505.38 192.49 510.01 ;
      RECT 191.69 35.31 192.29 35.51 ;
      RECT 191.77 30.13 192.09 30.73 ;
      RECT 191.77 42.75 192.09 43.35 ;
      RECT 183.69 28.15 191.89 28.75 ;
      RECT 191.09 59.37 191.73 59.97 ;
      RECT 172.79 35.75 191.69 35.95 ;
      RECT 172.79 37.21 191.69 37.41 ;
      RECT 191.49 63.99 191.69 505.18 ;
      RECT 191.49 505.38 191.69 510.01 ;
      RECT 172.79 34.65 191.49 34.85 ;
      RECT 191.09 505.38 191.29 510.01 ;
      RECT 189.21 6.24 191.19 6.84 ;
      RECT 190.49 35.31 191.09 35.51 ;
      RECT 190.69 30.13 191.01 30.73 ;
      RECT 190.69 42.75 191.01 43.35 ;
      RECT 190.29 505.38 190.49 510.01 ;
      RECT 189.89 505.38 190.09 510.01 ;
      RECT 189.29 35.31 189.89 35.51 ;
      RECT 189.37 30.13 189.69 30.73 ;
      RECT 189.37 42.75 189.69 43.35 ;
      RECT 189.49 65.96 189.69 510.01 ;
      RECT 188.65 59.37 189.29 59.97 ;
      RECT 189.09 505.38 189.29 510.01 ;
      RECT 188.69 63.99 188.89 505.18 ;
      RECT 188.69 505.38 188.89 510.01 ;
      RECT 186.81 6.24 188.79 6.84 ;
      RECT 188.09 35.31 188.69 35.51 ;
      RECT 188.29 30.13 188.61 30.73 ;
      RECT 188.29 42.75 188.61 43.35 ;
      RECT 187.09 15.51 188.49 15.71 ;
      RECT 188.29 65.96 188.49 510.01 ;
      RECT 187.89 505.38 188.09 510.01 ;
      RECT 187.49 505.38 187.69 510.01 ;
      RECT 186.89 35.31 187.49 35.51 ;
      RECT 186.97 30.13 187.29 30.73 ;
      RECT 186.97 42.75 187.29 43.35 ;
      RECT 186.29 59.37 186.93 59.97 ;
      RECT 186.69 63.99 186.89 505.18 ;
      RECT 186.69 505.38 186.89 510.01 ;
      RECT 186.29 505.38 186.49 510.01 ;
      RECT 184.41 6.24 186.39 6.84 ;
      RECT 185.69 35.31 186.29 35.51 ;
      RECT 185.89 30.13 186.21 30.73 ;
      RECT 185.89 42.75 186.21 43.35 ;
      RECT 185.49 505.38 185.69 510.01 ;
      RECT 185.09 505.38 185.29 510.01 ;
      RECT 184.49 35.31 185.09 35.51 ;
      RECT 184.57 30.13 184.89 30.73 ;
      RECT 184.57 42.75 184.89 43.35 ;
      RECT 184.69 65.96 184.89 510.01 ;
      RECT 183.85 59.37 184.49 59.97 ;
      RECT 184.29 505.38 184.49 510.01 ;
      RECT 183.89 63.99 184.09 505.18 ;
      RECT 183.89 505.38 184.09 510.01 ;
      RECT 181.99 6.24 183.99 6.84 ;
      RECT 183.29 35.31 183.89 35.51 ;
      RECT 183.49 30.13 183.81 30.73 ;
      RECT 183.49 42.75 183.81 43.35 ;
      RECT 183.49 65.96 183.69 510.01 ;
      RECT 182.83 12.98 183.43 13.18 ;
      RECT 183.09 505.38 183.29 510.01 ;
      RECT 182.69 505.38 182.89 510.01 ;
      RECT 181.73 8.94 182.69 9.14 ;
      RECT 182.09 35.31 182.69 35.51 ;
      RECT 178.23 13.78 182.59 13.98 ;
      RECT 182.17 30.13 182.49 30.73 ;
      RECT 182.17 42.75 182.49 43.35 ;
      RECT 182.14 28.03 182.34 28.77 ;
      RECT 174.19 21.31 182.19 21.51 ;
      RECT 180.23 20.61 182.18 21.01 ;
      RECT 181.49 59.37 182.13 59.97 ;
      RECT 181.89 63.99 182.09 505.18 ;
      RECT 181.89 505.38 182.09 510.01 ;
      RECT 180.9 16.58 181.94 16.78 ;
      RECT 174.44 27.51 181.94 27.71 ;
      RECT 174.44 27.91 181.94 28.11 ;
      RECT 181.49 505.38 181.69 510.01 ;
      RECT 179.62 6.24 181.59 6.84 ;
      RECT 180.89 35.31 181.49 35.51 ;
      RECT 174.91 22.31 181.47 22.51 ;
      RECT 181.09 30.13 181.41 30.73 ;
      RECT 181.09 42.75 181.41 43.35 ;
      RECT 175.15 9.98 181.27 10.18 ;
      RECT 180.15 23.11 181.19 23.31 ;
      RECT 173.89 13.38 181.07 13.58 ;
      RECT 180.29 28.72 180.89 28.92 ;
      RECT 180.69 505.38 180.89 510.01 ;
      RECT 180.15 8.94 180.75 9.14 ;
      RECT 180.29 505.38 180.49 510.01 ;
      RECT 179.38 15.39 180.46 15.59 ;
      RECT 176.03 28.31 180.35 28.51 ;
      RECT 179.69 35.31 180.29 35.51 ;
      RECT 179.59 12.98 180.19 13.18 ;
      RECT 179.77 30.13 180.09 30.73 ;
      RECT 179.77 42.75 180.09 43.35 ;
      RECT 179.89 65.96 180.09 510.01 ;
      RECT 179.73 24.3 179.93 25.07 ;
      RECT 176.53 20.79 179.85 20.99 ;
      RECT 179.05 59.37 179.69 59.97 ;
      RECT 179.49 505.38 179.69 510.01 ;
      RECT 177.59 8.94 179.31 9.14 ;
      RECT 179.09 63.99 179.29 505.18 ;
      RECT 179.09 505.38 179.29 510.01 ;
      RECT 177.69 6.24 179.19 6.84 ;
      RECT 178.49 35.31 179.09 35.51 ;
      RECT 178.69 30.13 179.01 30.73 ;
      RECT 178.69 42.75 179.01 43.35 ;
      RECT 178.69 65.96 178.89 510.01 ;
      RECT 177.79 15.38 178.79 15.72 ;
      RECT 177.63 20.38 178.75 20.58 ;
      RECT 178.29 505.38 178.49 510.01 ;
      RECT 177.89 505.38 178.09 510.01 ;
      RECT 177.29 35.31 177.89 35.51 ;
      RECT 177.37 30.13 177.69 30.73 ;
      RECT 177.37 42.75 177.69 43.35 ;
      RECT 173.79 16.5 177.65 16.7 ;
      RECT 175.79 15.38 177.47 15.58 ;
      RECT 176.79 8.94 177.39 9.14 ;
      RECT 176.69 59.37 177.33 59.97 ;
      RECT 177.09 63.99 177.29 505.18 ;
      RECT 177.09 505.38 177.29 510.01 ;
      RECT 176.69 505.38 176.89 510.01 ;
      RECT 175.27 12.58 176.69 12.78 ;
      RECT 176.09 35.31 176.69 35.51 ;
      RECT 176.45 24.3 176.65 25.07 ;
      RECT 176.29 30.13 176.61 30.73 ;
      RECT 176.29 42.75 176.61 43.35 ;
      RECT 175.79 18.61 176.39 18.81 ;
      RECT 175.29 6.24 176.29 6.84 ;
      RECT 175.19 23.11 176.23 23.31 ;
      RECT 174.2 20.61 176.15 21.01 ;
      RECT 175.49 28.72 176.09 28.92 ;
      RECT 175.89 505.38 176.09 510.01 ;
      RECT 175.49 505.38 175.69 510.01 ;
      RECT 174.89 35.31 175.49 35.51 ;
      RECT 174.97 30.13 175.29 30.73 ;
      RECT 174.97 42.75 175.29 43.35 ;
      RECT 175.09 65.96 175.29 510.01 ;
      RECT 174.25 59.37 174.89 59.97 ;
      RECT 174.69 505.38 174.89 510.01 ;
      RECT 174.29 63.99 174.49 505.18 ;
      RECT 174.29 505.38 174.49 510.01 ;
      RECT 173.69 35.31 174.29 35.51 ;
      RECT 174.04 28.03 174.24 28.77 ;
      RECT 173.89 30.13 174.21 30.73 ;
      RECT 173.89 42.75 174.21 43.35 ;
      RECT 173.89 65.96 174.09 510.01 ;
      RECT 173.79 15.38 173.99 15.98 ;
      RECT 172.99 6.24 173.79 6.84 ;
      RECT 173.49 505.38 173.69 510.01 ;
      RECT 173.29 12.58 173.49 13.85 ;
      RECT 173.09 505.38 173.29 510.01 ;
      RECT 172.49 35.31 173.09 35.51 ;
      RECT 172.79 15.38 172.99 15.98 ;
      RECT 169.13 16.5 172.99 16.7 ;
      RECT 165.71 13.38 172.89 13.58 ;
      RECT 172.57 30.13 172.89 30.73 ;
      RECT 172.57 42.75 172.89 43.35 ;
      RECT 172.54 28.03 172.74 28.77 ;
      RECT 164.59 21.31 172.59 21.51 ;
      RECT 170.63 20.61 172.58 21.01 ;
      RECT 171.89 59.37 172.53 59.97 ;
      RECT 154.19 35.75 172.49 35.95 ;
      RECT 154.19 37.21 172.49 37.41 ;
      RECT 172.29 63.99 172.49 505.18 ;
      RECT 172.29 505.38 172.49 510.01 ;
      RECT 164.84 27.51 172.34 27.71 ;
      RECT 164.84 27.91 172.34 28.11 ;
      RECT 154.19 34.65 172.29 34.85 ;
      RECT 171.89 505.38 172.09 510.01 ;
      RECT 171.29 35.31 171.89 35.51 ;
      RECT 165.31 22.31 171.87 22.51 ;
      RECT 171.49 30.13 171.81 30.73 ;
      RECT 171.49 42.75 171.81 43.35 ;
      RECT 165.51 9.98 171.63 10.18 ;
      RECT 170.55 23.11 171.59 23.31 ;
      RECT 170.09 12.58 171.51 12.78 ;
      RECT 170.49 6.24 171.49 6.84 ;
      RECT 170.69 28.72 171.29 28.92 ;
      RECT 171.09 505.38 171.29 510.01 ;
      RECT 169.31 15.38 170.99 15.58 ;
      RECT 170.39 18.61 170.99 18.81 ;
      RECT 170.69 505.38 170.89 510.01 ;
      RECT 166.43 28.31 170.75 28.51 ;
      RECT 170.09 35.31 170.69 35.51 ;
      RECT 170.17 30.13 170.49 30.73 ;
      RECT 170.17 42.75 170.49 43.35 ;
      RECT 170.29 65.96 170.49 510.01 ;
      RECT 170.13 24.3 170.33 25.07 ;
      RECT 166.93 20.79 170.25 20.99 ;
      RECT 169.45 59.37 170.09 59.97 ;
      RECT 169.89 505.38 170.09 510.01 ;
      RECT 169.39 8.94 169.99 9.14 ;
      RECT 169.49 63.99 169.69 505.18 ;
      RECT 169.49 505.38 169.69 510.01 ;
      RECT 168.89 35.31 169.49 35.51 ;
      RECT 169.09 30.13 169.41 30.73 ;
      RECT 169.09 42.75 169.41 43.35 ;
      RECT 169.09 65.96 169.29 510.01 ;
      RECT 167.47 8.94 169.19 9.14 ;
      RECT 168.03 20.38 169.15 20.58 ;
      RECT 167.59 6.24 169.09 6.84 ;
      RECT 167.99 15.38 168.99 15.72 ;
      RECT 168.69 505.38 168.89 510.01 ;
      RECT 164.19 13.78 168.55 13.98 ;
      RECT 168.29 505.38 168.49 510.01 ;
      RECT 167.69 35.31 168.29 35.51 ;
      RECT 167.77 30.13 168.09 30.73 ;
      RECT 167.77 42.75 168.09 43.35 ;
      RECT 167.09 59.37 167.73 59.97 ;
      RECT 167.49 63.99 167.69 505.18 ;
      RECT 167.49 505.38 167.69 510.01 ;
      RECT 166.32 15.39 167.4 15.59 ;
      RECT 167.09 505.38 167.29 510.01 ;
      RECT 166.59 12.98 167.19 13.18 ;
      RECT 165.19 6.24 167.16 6.84 ;
      RECT 166.49 35.31 167.09 35.51 ;
      RECT 166.85 24.3 167.05 25.07 ;
      RECT 166.69 30.13 167.01 30.73 ;
      RECT 166.69 42.75 167.01 43.35 ;
      RECT 166.03 8.94 166.63 9.14 ;
      RECT 165.59 23.11 166.63 23.31 ;
      RECT 164.6 20.61 166.55 21.01 ;
      RECT 165.89 28.72 166.49 28.92 ;
      RECT 166.29 505.38 166.49 510.01 ;
      RECT 165.89 505.38 166.09 510.01 ;
      RECT 165.29 35.31 165.89 35.51 ;
      RECT 164.84 16.58 165.88 16.78 ;
      RECT 165.37 30.13 165.69 30.73 ;
      RECT 165.37 42.75 165.69 43.35 ;
      RECT 165.49 65.96 165.69 510.01 ;
      RECT 164.65 59.37 165.29 59.97 ;
      RECT 165.09 505.38 165.29 510.01 ;
      RECT 164.09 8.94 165.05 9.14 ;
      RECT 164.69 63.99 164.89 505.18 ;
      RECT 164.69 505.38 164.89 510.01 ;
      RECT 162.79 6.24 164.79 6.84 ;
      RECT 164.09 35.31 164.69 35.51 ;
      RECT 164.44 28.03 164.64 28.77 ;
      RECT 164.29 30.13 164.61 30.73 ;
      RECT 164.29 42.75 164.61 43.35 ;
      RECT 164.29 65.96 164.49 510.01 ;
      RECT 163.89 505.38 164.09 510.01 ;
      RECT 163.35 12.98 163.95 13.18 ;
      RECT 163.49 505.38 163.69 510.01 ;
      RECT 162.89 35.31 163.49 35.51 ;
      RECT 162.97 30.13 163.29 30.73 ;
      RECT 162.97 42.75 163.29 43.35 ;
      RECT 154.89 28.15 163.09 28.75 ;
      RECT 162.29 59.37 162.93 59.97 ;
      RECT 162.69 63.99 162.89 505.18 ;
      RECT 162.69 505.38 162.89 510.01 ;
      RECT 162.29 505.38 162.49 510.01 ;
      RECT 160.39 6.24 162.37 6.84 ;
      RECT 161.69 35.31 162.29 35.51 ;
      RECT 161.89 30.13 162.21 30.73 ;
      RECT 161.89 42.75 162.21 43.35 ;
      RECT 161.49 505.38 161.69 510.01 ;
      RECT 161.09 505.38 161.29 510.01 ;
      RECT 160.49 35.31 161.09 35.51 ;
      RECT 160.57 30.13 160.89 30.73 ;
      RECT 160.57 42.75 160.89 43.35 ;
      RECT 160.69 65.96 160.89 510.01 ;
      RECT 159.85 59.37 160.49 59.97 ;
      RECT 160.29 505.38 160.49 510.01 ;
      RECT 159.89 63.99 160.09 505.18 ;
      RECT 159.89 505.38 160.09 510.01 ;
      RECT 157.99 6.24 159.97 6.84 ;
      RECT 159.29 35.31 159.89 35.51 ;
      RECT 159.49 30.13 159.81 30.73 ;
      RECT 159.49 42.75 159.81 43.35 ;
      RECT 158.29 15.51 159.69 15.71 ;
      RECT 159.49 65.96 159.69 510.01 ;
      RECT 159.09 505.38 159.29 510.01 ;
      RECT 158.69 505.38 158.89 510.01 ;
      RECT 158.09 35.31 158.69 35.51 ;
      RECT 158.17 30.13 158.49 30.73 ;
      RECT 158.17 42.75 158.49 43.35 ;
      RECT 157.49 59.37 158.13 59.97 ;
      RECT 157.89 63.99 158.09 505.18 ;
      RECT 157.89 505.38 158.09 510.01 ;
      RECT 157.49 505.38 157.69 510.01 ;
      RECT 155.59 6.24 157.57 6.84 ;
      RECT 156.89 35.31 157.49 35.51 ;
      RECT 157.09 30.13 157.41 30.73 ;
      RECT 157.09 42.75 157.41 43.35 ;
      RECT 156.69 505.38 156.89 510.01 ;
      RECT 156.29 505.38 156.49 510.01 ;
      RECT 155.69 35.31 156.29 35.51 ;
      RECT 155.77 30.13 156.09 30.73 ;
      RECT 155.77 42.75 156.09 43.35 ;
      RECT 155.89 65.96 156.09 510.01 ;
      RECT 155.05 59.37 155.69 59.97 ;
      RECT 155.49 505.38 155.69 510.01 ;
      RECT 155.09 63.99 155.29 505.18 ;
      RECT 155.09 505.38 155.29 510.01 ;
      RECT 153.89 6.24 155.19 6.84 ;
      RECT 154.49 35.31 155.09 35.51 ;
      RECT 154.69 30.13 155.01 30.73 ;
      RECT 154.69 42.75 155.01 43.35 ;
      RECT 154.69 65.96 154.89 510.01 ;
      RECT 154.29 505.38 154.49 510.01 ;
      RECT 153.49 68.06 153.69 70.14 ;
      RECT 153.49 70.34 153.69 71.16 ;
      RECT 153.49 71.36 153.69 72.18 ;
      RECT 153.49 72.38 153.69 73.54 ;
      RECT 153.49 73.74 153.69 74.56 ;
      RECT 153.49 74.76 153.69 75.58 ;
      RECT 153.49 75.78 153.69 76.94 ;
      RECT 153.49 77.14 153.69 77.96 ;
      RECT 153.49 78.16 153.69 78.98 ;
      RECT 153.49 79.18 153.69 80.34 ;
      RECT 153.49 80.54 153.69 81.36 ;
      RECT 153.49 81.56 153.69 82.38 ;
      RECT 153.49 82.58 153.69 83.74 ;
      RECT 153.49 83.94 153.69 84.76 ;
      RECT 153.49 84.96 153.69 85.78 ;
      RECT 153.49 85.98 153.69 87.14 ;
      RECT 153.49 87.34 153.69 88.16 ;
      RECT 153.49 88.36 153.69 89.18 ;
      RECT 153.49 89.38 153.69 90.54 ;
      RECT 153.49 90.74 153.69 91.56 ;
      RECT 153.49 91.76 153.69 92.58 ;
      RECT 153.49 92.78 153.69 93.94 ;
      RECT 153.49 94.14 153.69 94.96 ;
      RECT 153.49 95.16 153.69 95.98 ;
      RECT 153.49 96.18 153.69 97.34 ;
      RECT 153.49 97.54 153.69 98.36 ;
      RECT 153.49 98.56 153.69 99.38 ;
      RECT 153.49 99.58 153.69 100.74 ;
      RECT 153.49 100.94 153.69 101.76 ;
      RECT 153.49 101.96 153.69 102.78 ;
      RECT 153.49 102.98 153.69 104.14 ;
      RECT 153.49 104.34 153.69 105.16 ;
      RECT 153.49 105.36 153.69 106.18 ;
      RECT 153.49 106.38 153.69 107.54 ;
      RECT 153.49 107.74 153.69 108.56 ;
      RECT 153.49 108.76 153.69 109.58 ;
      RECT 153.49 109.78 153.69 110.94 ;
      RECT 153.49 111.14 153.69 111.96 ;
      RECT 153.49 112.16 153.69 112.98 ;
      RECT 153.49 113.18 153.69 114.34 ;
      RECT 153.49 114.54 153.69 115.36 ;
      RECT 153.49 115.56 153.69 116.38 ;
      RECT 153.49 116.58 153.69 117.74 ;
      RECT 153.49 117.94 153.69 118.76 ;
      RECT 153.49 118.96 153.69 119.78 ;
      RECT 153.49 119.98 153.69 121.14 ;
      RECT 153.49 121.34 153.69 122.16 ;
      RECT 153.49 122.36 153.69 123.18 ;
      RECT 153.49 123.38 153.69 124.54 ;
      RECT 153.49 124.74 153.69 125.56 ;
      RECT 153.49 125.76 153.69 126.58 ;
      RECT 153.49 126.78 153.69 127.94 ;
      RECT 153.49 128.14 153.69 128.96 ;
      RECT 153.49 129.16 153.69 129.98 ;
      RECT 153.49 130.18 153.69 131.34 ;
      RECT 153.49 131.54 153.69 132.36 ;
      RECT 153.49 132.56 153.69 133.38 ;
      RECT 153.49 133.58 153.69 134.74 ;
      RECT 153.49 134.94 153.69 135.76 ;
      RECT 153.49 135.96 153.69 136.78 ;
      RECT 153.49 136.98 153.69 138.14 ;
      RECT 153.49 138.34 153.69 139.16 ;
      RECT 153.49 139.36 153.69 140.18 ;
      RECT 153.49 140.38 153.69 141.54 ;
      RECT 153.49 141.74 153.69 142.56 ;
      RECT 153.49 142.76 153.69 143.58 ;
      RECT 153.49 143.78 153.69 144.94 ;
      RECT 153.49 145.14 153.69 145.96 ;
      RECT 153.49 146.16 153.69 146.98 ;
      RECT 153.49 147.18 153.69 148.34 ;
      RECT 153.49 148.54 153.69 149.36 ;
      RECT 153.49 149.56 153.69 150.38 ;
      RECT 153.49 150.58 153.69 151.74 ;
      RECT 153.49 151.94 153.69 152.76 ;
      RECT 153.49 152.96 153.69 153.78 ;
      RECT 153.49 153.98 153.69 155.14 ;
      RECT 153.49 155.34 153.69 156.16 ;
      RECT 153.49 156.36 153.69 157.18 ;
      RECT 153.49 157.38 153.69 158.54 ;
      RECT 153.49 158.74 153.69 159.56 ;
      RECT 153.49 159.76 153.69 160.58 ;
      RECT 153.49 160.78 153.69 161.94 ;
      RECT 153.49 162.14 153.69 162.96 ;
      RECT 153.49 163.16 153.69 163.98 ;
      RECT 153.49 164.18 153.69 165.34 ;
      RECT 153.49 165.54 153.69 166.36 ;
      RECT 153.49 166.56 153.69 167.38 ;
      RECT 153.49 167.58 153.69 168.74 ;
      RECT 153.49 168.94 153.69 169.76 ;
      RECT 153.49 169.96 153.69 170.78 ;
      RECT 153.49 170.98 153.69 172.14 ;
      RECT 153.49 172.34 153.69 173.16 ;
      RECT 153.49 173.36 153.69 174.18 ;
      RECT 153.49 174.38 153.69 175.54 ;
      RECT 153.49 175.74 153.69 176.56 ;
      RECT 153.49 176.76 153.69 177.58 ;
      RECT 153.49 177.78 153.69 178.94 ;
      RECT 153.49 179.14 153.69 179.96 ;
      RECT 153.49 180.16 153.69 180.98 ;
      RECT 153.49 181.18 153.69 182.34 ;
      RECT 153.49 182.54 153.69 183.36 ;
      RECT 153.49 183.56 153.69 184.38 ;
      RECT 153.49 184.58 153.69 185.74 ;
      RECT 153.49 185.94 153.69 186.76 ;
      RECT 153.49 186.96 153.69 187.78 ;
      RECT 153.49 187.98 153.69 189.14 ;
      RECT 153.49 189.34 153.69 190.16 ;
      RECT 153.49 190.36 153.69 191.18 ;
      RECT 153.49 191.38 153.69 192.54 ;
      RECT 153.49 192.74 153.69 193.56 ;
      RECT 153.49 193.76 153.69 194.58 ;
      RECT 153.49 194.78 153.69 195.94 ;
      RECT 153.49 196.14 153.69 196.96 ;
      RECT 153.49 197.16 153.69 197.98 ;
      RECT 153.49 198.18 153.69 199.34 ;
      RECT 153.49 199.54 153.69 200.36 ;
      RECT 153.49 200.56 153.69 201.38 ;
      RECT 153.49 201.58 153.69 202.74 ;
      RECT 153.49 202.94 153.69 203.76 ;
      RECT 153.49 203.96 153.69 204.78 ;
      RECT 153.49 204.98 153.69 206.14 ;
      RECT 153.49 206.34 153.69 207.16 ;
      RECT 153.49 207.36 153.69 208.18 ;
      RECT 153.49 208.38 153.69 209.54 ;
      RECT 153.49 209.74 153.69 210.56 ;
      RECT 153.49 210.76 153.69 211.58 ;
      RECT 153.49 211.78 153.69 212.94 ;
      RECT 153.49 213.14 153.69 213.96 ;
      RECT 153.49 214.16 153.69 214.98 ;
      RECT 153.49 215.18 153.69 216.34 ;
      RECT 153.49 216.54 153.69 217.36 ;
      RECT 153.49 217.56 153.69 218.38 ;
      RECT 153.49 218.58 153.69 219.74 ;
      RECT 153.49 219.94 153.69 220.76 ;
      RECT 153.49 220.96 153.69 221.78 ;
      RECT 153.49 221.98 153.69 223.14 ;
      RECT 153.49 223.34 153.69 224.16 ;
      RECT 153.49 224.36 153.69 225.18 ;
      RECT 153.49 225.38 153.69 226.54 ;
      RECT 153.49 226.74 153.69 227.56 ;
      RECT 153.49 227.76 153.69 228.58 ;
      RECT 153.49 228.78 153.69 229.94 ;
      RECT 153.49 230.14 153.69 230.96 ;
      RECT 153.49 231.16 153.69 231.98 ;
      RECT 153.49 232.18 153.69 233.34 ;
      RECT 153.49 233.54 153.69 234.36 ;
      RECT 153.49 234.56 153.69 235.38 ;
      RECT 153.49 235.58 153.69 236.74 ;
      RECT 153.49 236.94 153.69 237.76 ;
      RECT 153.49 237.96 153.69 238.78 ;
      RECT 153.49 238.98 153.69 240.14 ;
      RECT 153.49 240.34 153.69 241.16 ;
      RECT 153.49 241.36 153.69 242.18 ;
      RECT 153.49 242.38 153.69 243.54 ;
      RECT 153.49 243.74 153.69 244.56 ;
      RECT 153.49 244.76 153.69 245.58 ;
      RECT 153.49 245.78 153.69 246.94 ;
      RECT 153.49 247.14 153.69 247.96 ;
      RECT 153.49 248.16 153.69 248.98 ;
      RECT 153.49 249.18 153.69 250.34 ;
      RECT 153.49 250.54 153.69 251.36 ;
      RECT 153.49 251.56 153.69 252.38 ;
      RECT 153.49 252.58 153.69 253.74 ;
      RECT 153.49 253.94 153.69 254.76 ;
      RECT 153.49 254.96 153.69 255.78 ;
      RECT 153.49 255.98 153.69 257.14 ;
      RECT 153.49 257.34 153.69 258.16 ;
      RECT 153.49 258.36 153.69 259.18 ;
      RECT 153.49 259.38 153.69 260.54 ;
      RECT 153.49 260.74 153.69 261.56 ;
      RECT 153.49 261.76 153.69 262.58 ;
      RECT 153.49 262.78 153.69 263.94 ;
      RECT 153.49 264.14 153.69 264.96 ;
      RECT 153.49 265.16 153.69 265.98 ;
      RECT 153.49 266.18 153.69 267.34 ;
      RECT 153.49 267.54 153.69 268.36 ;
      RECT 153.49 268.56 153.69 269.38 ;
      RECT 153.49 269.58 153.69 270.74 ;
      RECT 153.49 270.94 153.69 271.76 ;
      RECT 153.49 271.96 153.69 272.78 ;
      RECT 153.49 272.98 153.69 274.14 ;
      RECT 153.49 274.34 153.69 275.16 ;
      RECT 153.49 275.36 153.69 276.18 ;
      RECT 153.49 276.38 153.69 277.54 ;
      RECT 153.49 277.74 153.69 278.56 ;
      RECT 153.49 278.76 153.69 279.58 ;
      RECT 153.49 279.78 153.69 280.94 ;
      RECT 153.49 281.14 153.69 281.96 ;
      RECT 153.49 282.16 153.69 282.98 ;
      RECT 153.49 283.18 153.69 284.34 ;
      RECT 153.49 284.54 153.69 285.36 ;
      RECT 153.49 285.56 153.69 286.38 ;
      RECT 153.49 286.58 153.69 287.74 ;
      RECT 153.49 287.94 153.69 288.76 ;
      RECT 153.49 288.96 153.69 289.78 ;
      RECT 153.49 289.98 153.69 291.14 ;
      RECT 153.49 291.34 153.69 292.16 ;
      RECT 153.49 292.36 153.69 293.18 ;
      RECT 153.49 293.38 153.69 294.54 ;
      RECT 153.49 294.74 153.69 295.56 ;
      RECT 153.49 295.76 153.69 296.58 ;
      RECT 153.49 296.78 153.69 297.94 ;
      RECT 153.49 298.14 153.69 298.96 ;
      RECT 153.49 299.16 153.69 299.98 ;
      RECT 153.49 300.18 153.69 301.34 ;
      RECT 153.49 301.54 153.69 302.36 ;
      RECT 153.49 302.56 153.69 303.38 ;
      RECT 153.49 303.58 153.69 304.74 ;
      RECT 153.49 304.94 153.69 305.76 ;
      RECT 153.49 305.96 153.69 306.78 ;
      RECT 153.49 306.98 153.69 308.14 ;
      RECT 153.49 308.34 153.69 309.16 ;
      RECT 153.49 309.36 153.69 310.18 ;
      RECT 153.49 310.38 153.69 311.54 ;
      RECT 153.49 311.74 153.69 312.56 ;
      RECT 153.49 312.76 153.69 313.58 ;
      RECT 153.49 313.78 153.69 314.94 ;
      RECT 153.49 315.14 153.69 315.96 ;
      RECT 153.49 316.16 153.69 316.98 ;
      RECT 153.49 317.18 153.69 318.34 ;
      RECT 153.49 318.54 153.69 319.36 ;
      RECT 153.49 319.56 153.69 320.38 ;
      RECT 153.49 320.58 153.69 321.74 ;
      RECT 153.49 321.94 153.69 322.76 ;
      RECT 153.49 322.96 153.69 323.78 ;
      RECT 153.49 323.98 153.69 325.14 ;
      RECT 153.49 325.34 153.69 326.16 ;
      RECT 153.49 326.36 153.69 327.18 ;
      RECT 153.49 327.38 153.69 328.54 ;
      RECT 153.49 328.74 153.69 329.56 ;
      RECT 153.49 329.76 153.69 330.58 ;
      RECT 153.49 330.78 153.69 331.94 ;
      RECT 153.49 332.14 153.69 332.96 ;
      RECT 153.49 333.16 153.69 333.98 ;
      RECT 153.49 334.18 153.69 335.34 ;
      RECT 153.49 335.54 153.69 336.36 ;
      RECT 153.49 336.56 153.69 337.38 ;
      RECT 153.49 337.58 153.69 338.74 ;
      RECT 153.49 338.94 153.69 339.76 ;
      RECT 153.49 339.96 153.69 340.78 ;
      RECT 153.49 340.98 153.69 342.14 ;
      RECT 153.49 342.34 153.69 343.16 ;
      RECT 153.49 343.36 153.69 344.18 ;
      RECT 153.49 344.38 153.69 345.54 ;
      RECT 153.49 345.74 153.69 346.56 ;
      RECT 153.49 346.76 153.69 347.58 ;
      RECT 153.49 347.78 153.69 348.94 ;
      RECT 153.49 349.14 153.69 349.96 ;
      RECT 153.49 350.16 153.69 350.98 ;
      RECT 153.49 351.18 153.69 352.34 ;
      RECT 153.49 352.54 153.69 353.36 ;
      RECT 153.49 353.56 153.69 354.38 ;
      RECT 153.49 354.58 153.69 355.74 ;
      RECT 153.49 355.94 153.69 356.76 ;
      RECT 153.49 356.96 153.69 357.78 ;
      RECT 153.49 357.98 153.69 359.14 ;
      RECT 153.49 359.34 153.69 360.16 ;
      RECT 153.49 360.36 153.69 361.18 ;
      RECT 153.49 361.38 153.69 362.54 ;
      RECT 153.49 362.74 153.69 363.56 ;
      RECT 153.49 363.76 153.69 364.58 ;
      RECT 153.49 364.78 153.69 365.94 ;
      RECT 153.49 366.14 153.69 366.96 ;
      RECT 153.49 367.16 153.69 367.98 ;
      RECT 153.49 368.18 153.69 369.34 ;
      RECT 153.49 369.54 153.69 370.36 ;
      RECT 153.49 370.56 153.69 371.38 ;
      RECT 153.49 371.58 153.69 372.74 ;
      RECT 153.49 372.94 153.69 373.76 ;
      RECT 153.49 373.96 153.69 374.78 ;
      RECT 153.49 374.98 153.69 376.14 ;
      RECT 153.49 376.34 153.69 377.16 ;
      RECT 153.49 377.36 153.69 378.18 ;
      RECT 153.49 378.38 153.69 379.54 ;
      RECT 153.49 379.74 153.69 380.56 ;
      RECT 153.49 380.76 153.69 381.58 ;
      RECT 153.49 381.78 153.69 382.94 ;
      RECT 153.49 383.14 153.69 383.96 ;
      RECT 153.49 384.16 153.69 384.98 ;
      RECT 153.49 385.18 153.69 386.34 ;
      RECT 153.49 386.54 153.69 387.36 ;
      RECT 153.49 387.56 153.69 388.38 ;
      RECT 153.49 388.58 153.69 389.74 ;
      RECT 153.49 389.94 153.69 390.76 ;
      RECT 153.49 390.96 153.69 391.78 ;
      RECT 153.49 391.98 153.69 393.14 ;
      RECT 153.49 393.34 153.69 394.16 ;
      RECT 153.49 394.36 153.69 395.18 ;
      RECT 153.49 395.38 153.69 396.54 ;
      RECT 153.49 396.74 153.69 397.56 ;
      RECT 153.49 397.76 153.69 398.58 ;
      RECT 153.49 398.78 153.69 399.94 ;
      RECT 153.49 400.14 153.69 400.96 ;
      RECT 153.49 401.16 153.69 401.98 ;
      RECT 153.49 402.18 153.69 403.34 ;
      RECT 153.49 403.54 153.69 404.36 ;
      RECT 153.49 404.56 153.69 405.38 ;
      RECT 153.49 405.58 153.69 406.74 ;
      RECT 153.49 406.94 153.69 407.76 ;
      RECT 153.49 407.96 153.69 408.78 ;
      RECT 153.49 408.98 153.69 410.14 ;
      RECT 153.49 410.34 153.69 411.16 ;
      RECT 153.49 411.36 153.69 412.18 ;
      RECT 153.49 412.38 153.69 413.54 ;
      RECT 153.49 413.74 153.69 414.56 ;
      RECT 153.49 414.76 153.69 415.58 ;
      RECT 153.49 415.78 153.69 416.94 ;
      RECT 153.49 417.14 153.69 417.96 ;
      RECT 153.49 418.16 153.69 418.98 ;
      RECT 153.49 419.18 153.69 420.34 ;
      RECT 153.49 420.54 153.69 421.36 ;
      RECT 153.49 421.56 153.69 422.38 ;
      RECT 153.49 422.58 153.69 423.74 ;
      RECT 153.49 423.94 153.69 424.76 ;
      RECT 153.49 424.96 153.69 425.78 ;
      RECT 153.49 425.98 153.69 427.14 ;
      RECT 153.49 427.34 153.69 428.16 ;
      RECT 153.49 428.36 153.69 429.18 ;
      RECT 153.49 429.38 153.69 430.54 ;
      RECT 153.49 430.74 153.69 431.56 ;
      RECT 153.49 431.76 153.69 432.58 ;
      RECT 153.49 432.78 153.69 433.94 ;
      RECT 153.49 434.14 153.69 434.96 ;
      RECT 153.49 435.16 153.69 435.98 ;
      RECT 153.49 436.18 153.69 437.34 ;
      RECT 153.49 437.54 153.69 438.36 ;
      RECT 153.49 438.56 153.69 439.38 ;
      RECT 153.49 439.58 153.69 440.74 ;
      RECT 153.49 440.94 153.69 441.76 ;
      RECT 153.49 441.96 153.69 442.78 ;
      RECT 153.49 442.98 153.69 444.14 ;
      RECT 153.49 444.34 153.69 445.16 ;
      RECT 153.49 445.36 153.69 446.18 ;
      RECT 153.49 446.38 153.69 447.54 ;
      RECT 153.49 447.74 153.69 448.56 ;
      RECT 153.49 448.76 153.69 449.58 ;
      RECT 153.49 449.78 153.69 450.94 ;
      RECT 153.49 451.14 153.69 451.96 ;
      RECT 153.49 452.16 153.69 452.98 ;
      RECT 153.49 453.18 153.69 454.34 ;
      RECT 153.49 454.54 153.69 455.36 ;
      RECT 153.49 455.56 153.69 456.38 ;
      RECT 153.49 456.58 153.69 457.74 ;
      RECT 153.49 457.94 153.69 458.76 ;
      RECT 153.49 458.96 153.69 459.78 ;
      RECT 153.49 459.98 153.69 461.14 ;
      RECT 153.49 461.34 153.69 462.16 ;
      RECT 153.49 462.36 153.69 463.18 ;
      RECT 153.49 463.38 153.69 464.54 ;
      RECT 153.49 464.74 153.69 465.56 ;
      RECT 153.49 465.76 153.69 466.58 ;
      RECT 153.49 466.78 153.69 467.94 ;
      RECT 153.49 468.14 153.69 468.96 ;
      RECT 153.49 469.16 153.69 469.98 ;
      RECT 153.49 470.18 153.69 471.34 ;
      RECT 153.49 471.54 153.69 472.36 ;
      RECT 153.49 472.56 153.69 473.38 ;
      RECT 153.49 473.58 153.69 474.74 ;
      RECT 153.49 474.94 153.69 475.76 ;
      RECT 153.49 475.96 153.69 476.78 ;
      RECT 153.49 476.98 153.69 478.14 ;
      RECT 153.49 478.34 153.69 479.16 ;
      RECT 153.49 479.36 153.69 480.18 ;
      RECT 153.49 480.38 153.69 481.54 ;
      RECT 153.49 481.74 153.69 482.56 ;
      RECT 153.49 482.76 153.69 483.58 ;
      RECT 153.49 483.78 153.69 484.94 ;
      RECT 153.49 485.14 153.69 485.96 ;
      RECT 153.49 486.16 153.69 486.98 ;
      RECT 153.49 487.18 153.69 488.34 ;
      RECT 153.49 488.54 153.69 489.36 ;
      RECT 153.49 489.56 153.69 490.38 ;
      RECT 153.49 490.58 153.69 491.74 ;
      RECT 153.49 491.94 153.69 492.76 ;
      RECT 153.49 492.96 153.69 493.78 ;
      RECT 153.49 493.98 153.69 495.14 ;
      RECT 153.49 495.34 153.69 496.16 ;
      RECT 153.49 496.36 153.69 497.18 ;
      RECT 153.49 497.38 153.69 498.54 ;
      RECT 153.49 498.74 153.69 499.56 ;
      RECT 153.49 499.76 153.69 500.58 ;
      RECT 153.49 500.78 153.69 501.94 ;
      RECT 153.49 502.14 153.69 502.96 ;
      RECT 153.49 503.16 153.69 503.98 ;
      RECT 153.49 504.18 153.69 506.38 ;
      RECT 153.49 506.58 153.69 507.4 ;
      RECT 153.49 507.6 153.69 508.42 ;
      RECT 153.49 508.62 153.69 510 ;
      RECT 152.89 23.74 153.49 23.94 ;
      RECT 149.18 16.27 153.41 16.47 ;
      RECT 152.57 22.64 153.15 22.92 ;
      RECT 140.49 42.85 153.09 43.15 ;
      RECT 152.69 68.06 152.89 510.06 ;
      RECT 151.99 510.34 152.79 510.94 ;
      RECT 148.59 29.95 152.69 30.15 ;
      RECT 152.29 68.06 152.49 507.66 ;
      RECT 140.49 43.54 152.31 43.84 ;
      RECT 149.89 16.96 152.11 17.16 ;
      RECT 151.89 68.06 152.09 509.06 ;
      RECT 141.97 23.71 151.93 24.74 ;
      RECT 145.99 32.44 151.91 32.64 ;
      RECT 151.29 6.24 151.89 6.84 ;
      RECT 147.98 27.51 151.89 27.71 ;
      RECT 140.39 51.67 151.79 51.87 ;
      RECT 151.49 68.06 151.69 507.66 ;
      RECT 145.17 22.86 151.62 23.06 ;
      RECT 150.79 510.34 151.59 510.94 ;
      RECT 88 31.15 151.54 32.15 ;
      RECT 150.71 22.39 151.49 22.59 ;
      RECT 150.85 30.75 151.49 30.95 ;
      RECT 88.21 63.23 151.47 65.03 ;
      RECT 151.09 68.06 151.29 70.14 ;
      RECT 151.09 70.34 151.29 72.18 ;
      RECT 151.09 72.38 151.29 73.54 ;
      RECT 151.09 73.74 151.29 75.58 ;
      RECT 151.09 75.78 151.29 76.94 ;
      RECT 151.09 77.14 151.29 78.98 ;
      RECT 151.09 79.18 151.29 80.34 ;
      RECT 151.09 80.54 151.29 82.38 ;
      RECT 151.09 82.58 151.29 83.74 ;
      RECT 151.09 83.94 151.29 85.78 ;
      RECT 151.09 85.98 151.29 87.14 ;
      RECT 151.09 87.34 151.29 89.18 ;
      RECT 151.09 89.38 151.29 90.54 ;
      RECT 151.09 90.74 151.29 92.58 ;
      RECT 151.09 92.78 151.29 93.94 ;
      RECT 151.09 94.14 151.29 95.98 ;
      RECT 151.09 96.18 151.29 97.34 ;
      RECT 151.09 97.54 151.29 99.38 ;
      RECT 151.09 99.58 151.29 100.74 ;
      RECT 151.09 100.94 151.29 102.78 ;
      RECT 151.09 102.98 151.29 104.14 ;
      RECT 151.09 104.34 151.29 106.18 ;
      RECT 151.09 106.38 151.29 107.54 ;
      RECT 151.09 107.74 151.29 109.58 ;
      RECT 151.09 109.78 151.29 110.94 ;
      RECT 151.09 111.14 151.29 112.98 ;
      RECT 151.09 113.18 151.29 114.34 ;
      RECT 151.09 114.54 151.29 116.38 ;
      RECT 151.09 116.58 151.29 117.74 ;
      RECT 151.09 117.94 151.29 119.78 ;
      RECT 151.09 119.98 151.29 121.14 ;
      RECT 151.09 121.34 151.29 123.18 ;
      RECT 151.09 123.38 151.29 124.54 ;
      RECT 151.09 124.74 151.29 126.58 ;
      RECT 151.09 126.78 151.29 127.94 ;
      RECT 151.09 128.14 151.29 129.98 ;
      RECT 151.09 130.18 151.29 131.34 ;
      RECT 151.09 131.54 151.29 133.38 ;
      RECT 151.09 133.58 151.29 134.74 ;
      RECT 151.09 134.94 151.29 136.78 ;
      RECT 151.09 136.98 151.29 138.14 ;
      RECT 151.09 138.34 151.29 140.18 ;
      RECT 151.09 140.38 151.29 141.54 ;
      RECT 151.09 141.74 151.29 143.58 ;
      RECT 151.09 143.78 151.29 144.94 ;
      RECT 151.09 145.14 151.29 146.98 ;
      RECT 151.09 147.18 151.29 148.34 ;
      RECT 151.09 148.54 151.29 150.38 ;
      RECT 151.09 150.58 151.29 151.74 ;
      RECT 151.09 151.94 151.29 153.78 ;
      RECT 151.09 153.98 151.29 155.14 ;
      RECT 151.09 155.34 151.29 157.18 ;
      RECT 151.09 157.38 151.29 158.54 ;
      RECT 151.09 158.74 151.29 160.58 ;
      RECT 151.09 160.78 151.29 161.94 ;
      RECT 151.09 162.14 151.29 163.98 ;
      RECT 151.09 164.18 151.29 165.34 ;
      RECT 151.09 165.54 151.29 167.38 ;
      RECT 151.09 167.58 151.29 168.74 ;
      RECT 151.09 168.94 151.29 170.78 ;
      RECT 151.09 170.98 151.29 172.14 ;
      RECT 151.09 172.34 151.29 174.18 ;
      RECT 151.09 174.38 151.29 175.54 ;
      RECT 151.09 175.74 151.29 177.58 ;
      RECT 151.09 177.78 151.29 178.94 ;
      RECT 151.09 179.14 151.29 180.98 ;
      RECT 151.09 181.18 151.29 182.34 ;
      RECT 151.09 182.54 151.29 184.38 ;
      RECT 151.09 184.58 151.29 185.74 ;
      RECT 151.09 185.94 151.29 187.78 ;
      RECT 151.09 187.98 151.29 189.14 ;
      RECT 151.09 189.34 151.29 191.18 ;
      RECT 151.09 191.38 151.29 192.54 ;
      RECT 151.09 192.74 151.29 194.58 ;
      RECT 151.09 194.78 151.29 195.94 ;
      RECT 151.09 196.14 151.29 197.98 ;
      RECT 151.09 198.18 151.29 199.34 ;
      RECT 151.09 199.54 151.29 201.38 ;
      RECT 151.09 201.58 151.29 202.74 ;
      RECT 151.09 202.94 151.29 204.78 ;
      RECT 151.09 204.98 151.29 206.14 ;
      RECT 151.09 206.34 151.29 208.18 ;
      RECT 151.09 208.38 151.29 209.54 ;
      RECT 151.09 209.74 151.29 211.58 ;
      RECT 151.09 211.78 151.29 212.94 ;
      RECT 151.09 213.14 151.29 214.98 ;
      RECT 151.09 215.18 151.29 216.34 ;
      RECT 151.09 216.54 151.29 218.38 ;
      RECT 151.09 218.58 151.29 219.74 ;
      RECT 151.09 219.94 151.29 221.78 ;
      RECT 151.09 221.98 151.29 223.14 ;
      RECT 151.09 223.34 151.29 225.18 ;
      RECT 151.09 225.38 151.29 226.54 ;
      RECT 151.09 226.74 151.29 228.58 ;
      RECT 151.09 228.78 151.29 229.94 ;
      RECT 151.09 230.14 151.29 231.98 ;
      RECT 151.09 232.18 151.29 233.34 ;
      RECT 151.09 233.54 151.29 235.38 ;
      RECT 151.09 235.58 151.29 236.74 ;
      RECT 151.09 236.94 151.29 238.78 ;
      RECT 151.09 238.98 151.29 240.14 ;
      RECT 151.09 240.34 151.29 242.18 ;
      RECT 151.09 242.38 151.29 243.54 ;
      RECT 151.09 243.74 151.29 245.58 ;
      RECT 151.09 245.78 151.29 246.94 ;
      RECT 151.09 247.14 151.29 248.98 ;
      RECT 151.09 249.18 151.29 250.34 ;
      RECT 151.09 250.54 151.29 252.38 ;
      RECT 151.09 252.58 151.29 253.74 ;
      RECT 151.09 253.94 151.29 255.78 ;
      RECT 151.09 255.98 151.29 257.14 ;
      RECT 151.09 257.34 151.29 259.18 ;
      RECT 151.09 259.38 151.29 260.54 ;
      RECT 151.09 260.74 151.29 262.58 ;
      RECT 151.09 262.78 151.29 263.94 ;
      RECT 151.09 264.14 151.29 265.98 ;
      RECT 151.09 266.18 151.29 267.34 ;
      RECT 151.09 267.54 151.29 269.38 ;
      RECT 151.09 269.58 151.29 270.74 ;
      RECT 151.09 270.94 151.29 272.78 ;
      RECT 151.09 272.98 151.29 274.14 ;
      RECT 151.09 274.34 151.29 276.18 ;
      RECT 151.09 276.38 151.29 277.54 ;
      RECT 151.09 277.74 151.29 279.58 ;
      RECT 151.09 279.78 151.29 280.94 ;
      RECT 151.09 281.14 151.29 282.98 ;
      RECT 151.09 283.18 151.29 284.34 ;
      RECT 151.09 284.54 151.29 286.38 ;
      RECT 151.09 286.58 151.29 287.74 ;
      RECT 151.09 287.94 151.29 289.78 ;
      RECT 151.09 289.98 151.29 291.14 ;
      RECT 151.09 291.34 151.29 293.18 ;
      RECT 151.09 293.38 151.29 294.54 ;
      RECT 151.09 294.74 151.29 296.58 ;
      RECT 151.09 296.78 151.29 297.94 ;
      RECT 151.09 298.14 151.29 299.98 ;
      RECT 151.09 300.18 151.29 301.34 ;
      RECT 151.09 301.54 151.29 303.38 ;
      RECT 151.09 303.58 151.29 304.74 ;
      RECT 151.09 304.94 151.29 306.78 ;
      RECT 151.09 306.98 151.29 308.14 ;
      RECT 151.09 308.34 151.29 310.18 ;
      RECT 151.09 310.38 151.29 311.54 ;
      RECT 151.09 311.74 151.29 313.58 ;
      RECT 151.09 313.78 151.29 314.94 ;
      RECT 151.09 315.14 151.29 316.98 ;
      RECT 151.09 317.18 151.29 318.34 ;
      RECT 151.09 318.54 151.29 320.38 ;
      RECT 151.09 320.58 151.29 321.74 ;
      RECT 151.09 321.94 151.29 323.78 ;
      RECT 151.09 323.98 151.29 325.14 ;
      RECT 151.09 325.34 151.29 327.18 ;
      RECT 151.09 327.38 151.29 328.54 ;
      RECT 151.09 328.74 151.29 330.58 ;
      RECT 151.09 330.78 151.29 331.94 ;
      RECT 151.09 332.14 151.29 333.98 ;
      RECT 151.09 334.18 151.29 335.34 ;
      RECT 151.09 335.54 151.29 337.38 ;
      RECT 151.09 337.58 151.29 338.74 ;
      RECT 151.09 338.94 151.29 340.78 ;
      RECT 151.09 340.98 151.29 342.14 ;
      RECT 151.09 342.34 151.29 344.18 ;
      RECT 151.09 344.38 151.29 345.54 ;
      RECT 151.09 345.74 151.29 347.58 ;
      RECT 151.09 347.78 151.29 348.94 ;
      RECT 151.09 349.14 151.29 350.98 ;
      RECT 151.09 351.18 151.29 352.34 ;
      RECT 151.09 352.54 151.29 354.38 ;
      RECT 151.09 354.58 151.29 355.74 ;
      RECT 151.09 355.94 151.29 357.78 ;
      RECT 151.09 357.98 151.29 359.14 ;
      RECT 151.09 359.34 151.29 361.18 ;
      RECT 151.09 361.38 151.29 362.54 ;
      RECT 151.09 362.74 151.29 364.58 ;
      RECT 151.09 364.78 151.29 365.94 ;
      RECT 151.09 366.14 151.29 367.98 ;
      RECT 151.09 368.18 151.29 369.34 ;
      RECT 151.09 369.54 151.29 371.38 ;
      RECT 151.09 371.58 151.29 372.74 ;
      RECT 151.09 372.94 151.29 374.78 ;
      RECT 151.09 374.98 151.29 376.14 ;
      RECT 151.09 376.34 151.29 378.18 ;
      RECT 151.09 378.38 151.29 379.54 ;
      RECT 151.09 379.74 151.29 381.58 ;
      RECT 151.09 381.78 151.29 382.94 ;
      RECT 151.09 383.14 151.29 384.98 ;
      RECT 151.09 385.18 151.29 386.34 ;
      RECT 151.09 386.54 151.29 388.38 ;
      RECT 151.09 388.58 151.29 389.74 ;
      RECT 151.09 389.94 151.29 391.78 ;
      RECT 151.09 391.98 151.29 393.14 ;
      RECT 151.09 393.34 151.29 395.18 ;
      RECT 151.09 395.38 151.29 396.54 ;
      RECT 151.09 396.74 151.29 398.58 ;
      RECT 151.09 398.78 151.29 399.94 ;
      RECT 151.09 400.14 151.29 401.98 ;
      RECT 151.09 402.18 151.29 403.34 ;
      RECT 151.09 403.54 151.29 405.38 ;
      RECT 151.09 405.58 151.29 406.74 ;
      RECT 151.09 406.94 151.29 408.78 ;
      RECT 151.09 408.98 151.29 410.14 ;
      RECT 151.09 410.34 151.29 412.18 ;
      RECT 151.09 412.38 151.29 413.54 ;
      RECT 151.09 413.74 151.29 415.58 ;
      RECT 151.09 415.78 151.29 416.94 ;
      RECT 151.09 417.14 151.29 418.98 ;
      RECT 151.09 419.18 151.29 420.34 ;
      RECT 151.09 420.54 151.29 422.38 ;
      RECT 151.09 422.58 151.29 423.74 ;
      RECT 151.09 423.94 151.29 425.78 ;
      RECT 151.09 425.98 151.29 427.14 ;
      RECT 151.09 427.34 151.29 429.18 ;
      RECT 151.09 429.38 151.29 430.54 ;
      RECT 151.09 430.74 151.29 432.58 ;
      RECT 151.09 432.78 151.29 433.94 ;
      RECT 151.09 434.14 151.29 435.98 ;
      RECT 151.09 436.18 151.29 437.34 ;
      RECT 151.09 437.54 151.29 439.38 ;
      RECT 151.09 439.58 151.29 440.74 ;
      RECT 151.09 440.94 151.29 442.78 ;
      RECT 151.09 442.98 151.29 444.14 ;
      RECT 151.09 444.34 151.29 446.18 ;
      RECT 151.09 446.38 151.29 447.54 ;
      RECT 151.09 447.74 151.29 449.58 ;
      RECT 151.09 449.78 151.29 450.94 ;
      RECT 151.09 451.14 151.29 452.98 ;
      RECT 151.09 453.18 151.29 454.34 ;
      RECT 151.09 454.54 151.29 456.38 ;
      RECT 151.09 456.58 151.29 457.74 ;
      RECT 151.09 457.94 151.29 459.78 ;
      RECT 151.09 459.98 151.29 461.14 ;
      RECT 151.09 461.34 151.29 463.18 ;
      RECT 151.09 463.38 151.29 464.54 ;
      RECT 151.09 464.74 151.29 466.58 ;
      RECT 151.09 466.78 151.29 467.94 ;
      RECT 151.09 468.14 151.29 469.98 ;
      RECT 151.09 470.18 151.29 471.34 ;
      RECT 151.09 471.54 151.29 473.38 ;
      RECT 151.09 473.58 151.29 474.74 ;
      RECT 151.09 474.94 151.29 476.78 ;
      RECT 151.09 476.98 151.29 478.14 ;
      RECT 151.09 478.34 151.29 480.18 ;
      RECT 151.09 480.38 151.29 481.54 ;
      RECT 151.09 481.74 151.29 483.58 ;
      RECT 151.09 483.78 151.29 484.94 ;
      RECT 151.09 485.14 151.29 486.98 ;
      RECT 151.09 487.18 151.29 488.34 ;
      RECT 151.09 488.54 151.29 490.38 ;
      RECT 151.09 490.58 151.29 491.74 ;
      RECT 151.09 491.94 151.29 493.78 ;
      RECT 151.09 493.98 151.29 495.14 ;
      RECT 151.09 495.34 151.29 497.18 ;
      RECT 151.09 497.38 151.29 498.54 ;
      RECT 151.09 498.74 151.29 500.58 ;
      RECT 151.09 500.78 151.29 501.94 ;
      RECT 151.09 502.14 151.29 503.98 ;
      RECT 151.09 504.18 151.29 505.96 ;
      RECT 140.39 35.34 151.19 35.54 ;
      RECT 147.65 29.46 151.11 29.66 ;
      RECT 143.81 25.43 151.09 25.63 ;
      RECT 150.29 6.24 150.89 6.84 ;
      RECT 150.69 68.06 150.89 507.66 ;
      RECT 109.39 68.83 150.49 69.03 ;
      RECT 150.16 69.41 150.42 69.96 ;
      RECT 150.16 72.56 150.42 73.36 ;
      RECT 150.16 75.96 150.42 76.76 ;
      RECT 150.16 79.36 150.42 80.16 ;
      RECT 150.16 82.76 150.42 83.56 ;
      RECT 150.16 86.16 150.42 86.96 ;
      RECT 150.16 89.56 150.42 90.36 ;
      RECT 150.16 92.96 150.42 93.76 ;
      RECT 150.16 96.36 150.42 97.16 ;
      RECT 150.16 99.76 150.42 100.56 ;
      RECT 150.16 103.16 150.42 103.96 ;
      RECT 150.16 106.56 150.42 107.36 ;
      RECT 150.16 109.96 150.42 110.76 ;
      RECT 150.16 113.36 150.42 114.16 ;
      RECT 150.16 116.76 150.42 117.56 ;
      RECT 150.16 120.16 150.42 120.96 ;
      RECT 150.16 123.56 150.42 124.36 ;
      RECT 150.16 126.96 150.42 127.76 ;
      RECT 150.16 130.36 150.42 131.16 ;
      RECT 150.16 133.76 150.42 134.56 ;
      RECT 150.16 137.16 150.42 137.96 ;
      RECT 150.16 140.56 150.42 141.36 ;
      RECT 150.16 143.96 150.42 144.76 ;
      RECT 150.16 147.36 150.42 148.16 ;
      RECT 150.16 150.76 150.42 151.56 ;
      RECT 150.16 154.16 150.42 154.96 ;
      RECT 150.16 157.56 150.42 158.36 ;
      RECT 150.16 160.96 150.42 161.76 ;
      RECT 150.16 164.36 150.42 165.16 ;
      RECT 150.16 167.76 150.42 168.56 ;
      RECT 150.16 171.16 150.42 171.96 ;
      RECT 150.16 174.56 150.42 175.36 ;
      RECT 150.16 177.96 150.42 178.76 ;
      RECT 150.16 181.36 150.42 182.16 ;
      RECT 150.16 184.76 150.42 185.56 ;
      RECT 150.16 188.16 150.42 188.96 ;
      RECT 150.16 191.56 150.42 192.36 ;
      RECT 150.16 194.96 150.42 195.76 ;
      RECT 150.16 198.36 150.42 199.16 ;
      RECT 150.16 201.76 150.42 202.56 ;
      RECT 150.16 205.16 150.42 205.96 ;
      RECT 150.16 208.56 150.42 209.36 ;
      RECT 150.16 211.96 150.42 212.76 ;
      RECT 150.16 215.36 150.42 216.16 ;
      RECT 150.16 218.76 150.42 219.56 ;
      RECT 150.16 222.16 150.42 222.96 ;
      RECT 150.16 225.56 150.42 226.36 ;
      RECT 150.16 228.96 150.42 229.76 ;
      RECT 150.16 232.36 150.42 233.16 ;
      RECT 150.16 235.76 150.42 236.56 ;
      RECT 150.16 239.16 150.42 239.96 ;
      RECT 150.16 242.56 150.42 243.36 ;
      RECT 150.16 245.96 150.42 246.76 ;
      RECT 150.16 249.36 150.42 250.16 ;
      RECT 150.16 252.76 150.42 253.56 ;
      RECT 150.16 256.16 150.42 256.96 ;
      RECT 150.16 259.56 150.42 260.36 ;
      RECT 150.16 262.96 150.42 263.76 ;
      RECT 150.16 266.36 150.42 267.16 ;
      RECT 150.16 269.76 150.42 270.56 ;
      RECT 150.16 273.16 150.42 273.96 ;
      RECT 150.16 276.56 150.42 277.36 ;
      RECT 150.16 279.96 150.42 280.76 ;
      RECT 150.16 283.36 150.42 284.16 ;
      RECT 150.16 286.76 150.42 287.56 ;
      RECT 150.16 290.16 150.42 290.96 ;
      RECT 150.16 293.56 150.42 294.36 ;
      RECT 150.16 296.96 150.42 297.76 ;
      RECT 150.16 300.36 150.42 301.16 ;
      RECT 150.16 303.76 150.42 304.56 ;
      RECT 150.16 307.16 150.42 307.96 ;
      RECT 150.16 310.56 150.42 311.36 ;
      RECT 150.16 313.96 150.42 314.76 ;
      RECT 150.16 317.36 150.42 318.16 ;
      RECT 150.16 320.76 150.42 321.56 ;
      RECT 150.16 324.16 150.42 324.96 ;
      RECT 150.16 327.56 150.42 328.36 ;
      RECT 150.16 330.96 150.42 331.76 ;
      RECT 150.16 334.36 150.42 335.16 ;
      RECT 150.16 337.76 150.42 338.56 ;
      RECT 150.16 341.16 150.42 341.96 ;
      RECT 150.16 344.56 150.42 345.36 ;
      RECT 150.16 347.96 150.42 348.76 ;
      RECT 150.16 351.36 150.42 352.16 ;
      RECT 150.16 354.76 150.42 355.56 ;
      RECT 150.16 358.16 150.42 358.96 ;
      RECT 150.16 361.56 150.42 362.36 ;
      RECT 150.16 364.96 150.42 365.76 ;
      RECT 150.16 368.36 150.42 369.16 ;
      RECT 150.16 371.76 150.42 372.56 ;
      RECT 150.16 375.16 150.42 375.96 ;
      RECT 150.16 378.56 150.42 379.36 ;
      RECT 150.16 381.96 150.42 382.76 ;
      RECT 150.16 385.36 150.42 386.16 ;
      RECT 150.16 388.76 150.42 389.56 ;
      RECT 150.16 392.16 150.42 392.96 ;
      RECT 150.16 395.56 150.42 396.36 ;
      RECT 150.16 398.96 150.42 399.76 ;
      RECT 150.16 402.36 150.42 403.16 ;
      RECT 150.16 405.76 150.42 406.56 ;
      RECT 150.16 409.16 150.42 409.96 ;
      RECT 150.16 412.56 150.42 413.36 ;
      RECT 150.16 415.96 150.42 416.76 ;
      RECT 150.16 419.36 150.42 420.16 ;
      RECT 150.16 422.76 150.42 423.56 ;
      RECT 150.16 426.16 150.42 426.96 ;
      RECT 150.16 429.56 150.42 430.36 ;
      RECT 150.16 432.96 150.42 433.76 ;
      RECT 150.16 436.36 150.42 437.16 ;
      RECT 150.16 439.76 150.42 440.56 ;
      RECT 150.16 443.16 150.42 443.96 ;
      RECT 150.16 446.56 150.42 447.36 ;
      RECT 150.16 449.96 150.42 450.76 ;
      RECT 150.16 453.36 150.42 454.16 ;
      RECT 150.16 456.76 150.42 457.56 ;
      RECT 150.16 460.16 150.42 460.96 ;
      RECT 150.16 463.56 150.42 464.36 ;
      RECT 150.16 466.96 150.42 467.76 ;
      RECT 150.16 470.36 150.42 471.16 ;
      RECT 150.16 473.76 150.42 474.56 ;
      RECT 150.16 477.16 150.42 477.96 ;
      RECT 150.16 480.56 150.42 481.36 ;
      RECT 150.16 483.96 150.42 484.76 ;
      RECT 150.16 487.36 150.42 488.16 ;
      RECT 150.16 490.76 150.42 491.56 ;
      RECT 150.16 494.16 150.42 494.96 ;
      RECT 150.16 497.56 150.42 498.36 ;
      RECT 150.16 500.96 150.42 501.76 ;
      RECT 150.16 504.36 150.42 504.91 ;
      RECT 149.66 70.96 150.41 71.56 ;
      RECT 149.66 74.36 150.41 74.96 ;
      RECT 149.66 77.76 150.41 78.36 ;
      RECT 149.66 81.16 150.41 81.76 ;
      RECT 149.66 84.56 150.41 85.16 ;
      RECT 149.66 87.96 150.41 88.56 ;
      RECT 149.66 91.36 150.41 91.96 ;
      RECT 149.66 94.76 150.41 95.36 ;
      RECT 149.66 98.16 150.41 98.76 ;
      RECT 149.66 101.56 150.41 102.16 ;
      RECT 149.66 104.96 150.41 105.56 ;
      RECT 149.66 108.36 150.41 108.96 ;
      RECT 149.66 111.76 150.41 112.36 ;
      RECT 149.66 115.16 150.41 115.76 ;
      RECT 149.66 118.56 150.41 119.16 ;
      RECT 149.66 121.96 150.41 122.56 ;
      RECT 149.66 125.36 150.41 125.96 ;
      RECT 149.66 128.76 150.41 129.36 ;
      RECT 149.66 132.16 150.41 132.76 ;
      RECT 149.66 135.56 150.41 136.16 ;
      RECT 149.66 138.96 150.41 139.56 ;
      RECT 149.66 142.36 150.41 142.96 ;
      RECT 149.66 145.76 150.41 146.36 ;
      RECT 149.66 149.16 150.41 149.76 ;
      RECT 149.66 152.56 150.41 153.16 ;
      RECT 149.66 155.96 150.41 156.56 ;
      RECT 149.66 159.36 150.41 159.96 ;
      RECT 149.66 162.76 150.41 163.36 ;
      RECT 149.66 166.16 150.41 166.76 ;
      RECT 149.66 169.56 150.41 170.16 ;
      RECT 149.66 172.96 150.41 173.56 ;
      RECT 149.66 176.36 150.41 176.96 ;
      RECT 149.66 179.76 150.41 180.36 ;
      RECT 149.66 183.16 150.41 183.76 ;
      RECT 149.66 186.56 150.41 187.16 ;
      RECT 149.66 189.96 150.41 190.56 ;
      RECT 149.66 193.36 150.41 193.96 ;
      RECT 149.66 196.76 150.41 197.36 ;
      RECT 149.66 200.16 150.41 200.76 ;
      RECT 149.66 203.56 150.41 204.16 ;
      RECT 149.66 206.96 150.41 207.56 ;
      RECT 149.66 210.36 150.41 210.96 ;
      RECT 149.66 213.76 150.41 214.36 ;
      RECT 149.66 217.16 150.41 217.76 ;
      RECT 149.66 220.56 150.41 221.16 ;
      RECT 149.66 223.96 150.41 224.56 ;
      RECT 149.66 227.36 150.41 227.96 ;
      RECT 149.66 230.76 150.41 231.36 ;
      RECT 149.66 234.16 150.41 234.76 ;
      RECT 149.66 237.56 150.41 238.16 ;
      RECT 149.66 240.96 150.41 241.56 ;
      RECT 149.66 244.36 150.41 244.96 ;
      RECT 149.66 247.76 150.41 248.36 ;
      RECT 149.66 251.16 150.41 251.76 ;
      RECT 149.66 254.56 150.41 255.16 ;
      RECT 149.66 257.96 150.41 258.56 ;
      RECT 149.66 261.36 150.41 261.96 ;
      RECT 149.66 264.76 150.41 265.36 ;
      RECT 149.66 268.16 150.41 268.76 ;
      RECT 149.66 271.56 150.41 272.16 ;
      RECT 149.66 274.96 150.41 275.56 ;
      RECT 149.66 278.36 150.41 278.96 ;
      RECT 149.66 281.76 150.41 282.36 ;
      RECT 149.66 285.16 150.41 285.76 ;
      RECT 149.66 288.56 150.41 289.16 ;
      RECT 149.66 291.96 150.41 292.56 ;
      RECT 149.66 295.36 150.41 295.96 ;
      RECT 149.66 298.76 150.41 299.36 ;
      RECT 149.66 302.16 150.41 302.76 ;
      RECT 149.66 305.56 150.41 306.16 ;
      RECT 149.66 308.96 150.41 309.56 ;
      RECT 149.66 312.36 150.41 312.96 ;
      RECT 149.66 315.76 150.41 316.36 ;
      RECT 149.66 319.16 150.41 319.76 ;
      RECT 149.66 322.56 150.41 323.16 ;
      RECT 149.66 325.96 150.41 326.56 ;
      RECT 149.66 329.36 150.41 329.96 ;
      RECT 149.66 332.76 150.41 333.36 ;
      RECT 149.66 336.16 150.41 336.76 ;
      RECT 149.66 339.56 150.41 340.16 ;
      RECT 149.66 342.96 150.41 343.56 ;
      RECT 149.66 346.36 150.41 346.96 ;
      RECT 149.66 349.76 150.41 350.36 ;
      RECT 149.66 353.16 150.41 353.76 ;
      RECT 149.66 356.56 150.41 357.16 ;
      RECT 149.66 359.96 150.41 360.56 ;
      RECT 149.66 363.36 150.41 363.96 ;
      RECT 149.66 366.76 150.41 367.36 ;
      RECT 149.66 370.16 150.41 370.76 ;
      RECT 149.66 373.56 150.41 374.16 ;
      RECT 149.66 376.96 150.41 377.56 ;
      RECT 149.66 380.36 150.41 380.96 ;
      RECT 149.66 383.76 150.41 384.36 ;
      RECT 149.66 387.16 150.41 387.76 ;
      RECT 149.66 390.56 150.41 391.16 ;
      RECT 149.66 393.96 150.41 394.56 ;
      RECT 149.66 397.36 150.41 397.96 ;
      RECT 149.66 400.76 150.41 401.36 ;
      RECT 149.66 404.16 150.41 404.76 ;
      RECT 149.66 407.56 150.41 408.16 ;
      RECT 149.66 410.96 150.41 411.56 ;
      RECT 149.66 414.36 150.41 414.96 ;
      RECT 149.66 417.76 150.41 418.36 ;
      RECT 149.66 421.16 150.41 421.76 ;
      RECT 149.66 424.56 150.41 425.16 ;
      RECT 149.66 427.96 150.41 428.56 ;
      RECT 149.66 431.36 150.41 431.96 ;
      RECT 149.66 434.76 150.41 435.36 ;
      RECT 149.66 438.16 150.41 438.76 ;
      RECT 149.66 441.56 150.41 442.16 ;
      RECT 149.66 444.96 150.41 445.56 ;
      RECT 149.66 448.36 150.41 448.96 ;
      RECT 149.66 451.76 150.41 452.36 ;
      RECT 149.66 455.16 150.41 455.76 ;
      RECT 149.66 458.56 150.41 459.16 ;
      RECT 149.66 461.96 150.41 462.56 ;
      RECT 149.66 465.36 150.41 465.96 ;
      RECT 149.66 468.76 150.41 469.36 ;
      RECT 149.66 472.16 150.41 472.76 ;
      RECT 149.66 475.56 150.41 476.16 ;
      RECT 149.66 478.96 150.41 479.56 ;
      RECT 149.66 482.36 150.41 482.96 ;
      RECT 149.66 485.76 150.41 486.36 ;
      RECT 149.66 489.16 150.41 489.76 ;
      RECT 149.66 492.56 150.41 493.16 ;
      RECT 149.66 495.96 150.41 496.56 ;
      RECT 149.66 499.36 150.41 499.96 ;
      RECT 149.66 502.76 150.41 503.36 ;
      RECT 149.93 510.34 150.39 510.94 ;
      RECT 148.9 52.16 150.38 52.76 ;
      RECT 145.65 30.75 150.05 30.95 ;
      RECT 149.43 508.1 149.85 508.6 ;
      RECT 149.49 62.18 149.77 62.78 ;
      RECT 145.65 27.91 149.39 28.11 ;
      RECT 148.01 510.34 149.33 510.94 ;
      RECT 148.05 10.23 149.29 10.83 ;
      RECT 131.61 69.46 149.29 69.66 ;
      RECT 131.61 72.86 149.29 73.06 ;
      RECT 131.61 76.26 149.29 76.46 ;
      RECT 131.61 79.66 149.29 79.86 ;
      RECT 131.61 83.06 149.29 83.26 ;
      RECT 131.61 86.46 149.29 86.66 ;
      RECT 131.61 89.86 149.29 90.06 ;
      RECT 131.61 93.26 149.29 93.46 ;
      RECT 131.61 96.66 149.29 96.86 ;
      RECT 131.61 100.06 149.29 100.26 ;
      RECT 131.61 103.46 149.29 103.66 ;
      RECT 131.61 106.86 149.29 107.06 ;
      RECT 131.61 110.26 149.29 110.46 ;
      RECT 131.61 113.66 149.29 113.86 ;
      RECT 131.61 117.06 149.29 117.26 ;
      RECT 131.61 120.46 149.29 120.66 ;
      RECT 131.61 123.86 149.29 124.06 ;
      RECT 131.61 127.26 149.29 127.46 ;
      RECT 131.61 130.66 149.29 130.86 ;
      RECT 131.61 134.06 149.29 134.26 ;
      RECT 131.61 137.46 149.29 137.66 ;
      RECT 131.61 140.86 149.29 141.06 ;
      RECT 131.61 144.26 149.29 144.46 ;
      RECT 131.61 147.66 149.29 147.86 ;
      RECT 131.61 151.06 149.29 151.26 ;
      RECT 131.61 154.46 149.29 154.66 ;
      RECT 131.61 157.86 149.29 158.06 ;
      RECT 131.61 161.26 149.29 161.46 ;
      RECT 131.61 164.66 149.29 164.86 ;
      RECT 131.61 168.06 149.29 168.26 ;
      RECT 131.61 171.46 149.29 171.66 ;
      RECT 131.61 174.86 149.29 175.06 ;
      RECT 131.61 178.26 149.29 178.46 ;
      RECT 131.61 181.66 149.29 181.86 ;
      RECT 131.61 185.06 149.29 185.26 ;
      RECT 131.61 188.46 149.29 188.66 ;
      RECT 131.61 191.86 149.29 192.06 ;
      RECT 131.61 195.26 149.29 195.46 ;
      RECT 131.61 198.66 149.29 198.86 ;
      RECT 131.61 202.06 149.29 202.26 ;
      RECT 131.61 205.46 149.29 205.66 ;
      RECT 131.61 208.86 149.29 209.06 ;
      RECT 131.61 212.26 149.29 212.46 ;
      RECT 131.61 215.66 149.29 215.86 ;
      RECT 131.61 219.06 149.29 219.26 ;
      RECT 131.61 222.46 149.29 222.66 ;
      RECT 131.61 225.86 149.29 226.06 ;
      RECT 131.61 229.26 149.29 229.46 ;
      RECT 131.61 232.66 149.29 232.86 ;
      RECT 131.61 236.06 149.29 236.26 ;
      RECT 131.61 239.46 149.29 239.66 ;
      RECT 131.61 242.86 149.29 243.06 ;
      RECT 131.61 246.26 149.29 246.46 ;
      RECT 131.61 249.66 149.29 249.86 ;
      RECT 131.61 253.06 149.29 253.26 ;
      RECT 131.61 256.46 149.29 256.66 ;
      RECT 131.61 259.86 149.29 260.06 ;
      RECT 131.61 263.26 149.29 263.46 ;
      RECT 131.61 266.66 149.29 266.86 ;
      RECT 131.61 270.06 149.29 270.26 ;
      RECT 131.61 273.46 149.29 273.66 ;
      RECT 131.61 276.86 149.29 277.06 ;
      RECT 131.61 280.26 149.29 280.46 ;
      RECT 131.61 283.66 149.29 283.86 ;
      RECT 131.61 287.06 149.29 287.26 ;
      RECT 131.61 290.46 149.29 290.66 ;
      RECT 131.61 293.86 149.29 294.06 ;
      RECT 131.61 297.26 149.29 297.46 ;
      RECT 131.61 300.66 149.29 300.86 ;
      RECT 131.61 304.06 149.29 304.26 ;
      RECT 131.61 307.46 149.29 307.66 ;
      RECT 131.61 310.86 149.29 311.06 ;
      RECT 131.61 314.26 149.29 314.46 ;
      RECT 131.61 317.66 149.29 317.86 ;
      RECT 131.61 321.06 149.29 321.26 ;
      RECT 131.61 324.46 149.29 324.66 ;
      RECT 131.61 327.86 149.29 328.06 ;
      RECT 131.61 331.26 149.29 331.46 ;
      RECT 131.61 334.66 149.29 334.86 ;
      RECT 131.61 338.06 149.29 338.26 ;
      RECT 131.61 341.46 149.29 341.66 ;
      RECT 131.61 344.86 149.29 345.06 ;
      RECT 131.61 348.26 149.29 348.46 ;
      RECT 131.61 351.66 149.29 351.86 ;
      RECT 131.61 355.06 149.29 355.26 ;
      RECT 131.61 358.46 149.29 358.66 ;
      RECT 131.61 361.86 149.29 362.06 ;
      RECT 131.61 365.26 149.29 365.46 ;
      RECT 131.61 368.66 149.29 368.86 ;
      RECT 131.61 372.06 149.29 372.26 ;
      RECT 131.61 375.46 149.29 375.66 ;
      RECT 131.61 378.86 149.29 379.06 ;
      RECT 131.61 382.26 149.29 382.46 ;
      RECT 131.61 385.66 149.29 385.86 ;
      RECT 131.61 389.06 149.29 389.26 ;
      RECT 131.61 392.46 149.29 392.66 ;
      RECT 131.61 395.86 149.29 396.06 ;
      RECT 131.61 399.26 149.29 399.46 ;
      RECT 131.61 402.66 149.29 402.86 ;
      RECT 131.61 406.06 149.29 406.26 ;
      RECT 131.61 409.46 149.29 409.66 ;
      RECT 131.61 412.86 149.29 413.06 ;
      RECT 131.61 416.26 149.29 416.46 ;
      RECT 131.61 419.66 149.29 419.86 ;
      RECT 131.61 423.06 149.29 423.26 ;
      RECT 131.61 426.46 149.29 426.66 ;
      RECT 131.61 429.86 149.29 430.06 ;
      RECT 131.61 433.26 149.29 433.46 ;
      RECT 131.61 436.66 149.29 436.86 ;
      RECT 131.61 440.06 149.29 440.26 ;
      RECT 131.61 443.46 149.29 443.66 ;
      RECT 131.61 446.86 149.29 447.06 ;
      RECT 131.61 450.26 149.29 450.46 ;
      RECT 131.61 453.66 149.29 453.86 ;
      RECT 131.61 457.06 149.29 457.26 ;
      RECT 131.61 460.46 149.29 460.66 ;
      RECT 131.61 463.86 149.29 464.06 ;
      RECT 131.61 467.26 149.29 467.46 ;
      RECT 131.61 470.66 149.29 470.86 ;
      RECT 131.61 474.06 149.29 474.26 ;
      RECT 131.61 477.46 149.29 477.66 ;
      RECT 131.61 480.86 149.29 481.06 ;
      RECT 131.61 484.26 149.29 484.46 ;
      RECT 131.61 487.66 149.29 487.86 ;
      RECT 131.61 491.06 149.29 491.26 ;
      RECT 131.61 494.46 149.29 494.66 ;
      RECT 131.61 497.86 149.29 498.06 ;
      RECT 131.61 501.26 149.29 501.46 ;
      RECT 131.61 504.66 149.29 504.86 ;
      RECT 137.99 506.86 149.01 507.38 ;
      RECT 148.01 6.24 148.87 6.84 ;
      RECT 135.41 508.7 148.81 509.22 ;
      RECT 137.99 509.42 148.81 509.94 ;
      RECT 146.96 52.16 148.44 52.76 ;
      RECT 146.06 16.27 147.85 16.47 ;
      RECT 147.57 62.18 147.85 62.78 ;
      RECT 146.09 6.24 147.41 6.84 ;
      RECT 146.09 70.42 147.41 70.62 ;
      RECT 146.09 71.9 147.41 72.1 ;
      RECT 146.09 73.82 147.41 74.02 ;
      RECT 146.09 75.3 147.41 75.5 ;
      RECT 146.09 77.22 147.41 77.42 ;
      RECT 146.09 78.7 147.41 78.9 ;
      RECT 146.09 80.62 147.41 80.82 ;
      RECT 146.09 82.1 147.41 82.3 ;
      RECT 146.09 84.02 147.41 84.22 ;
      RECT 146.09 85.5 147.41 85.7 ;
      RECT 146.09 87.42 147.41 87.62 ;
      RECT 146.09 88.9 147.41 89.1 ;
      RECT 146.09 90.82 147.41 91.02 ;
      RECT 146.09 92.3 147.41 92.5 ;
      RECT 146.09 94.22 147.41 94.42 ;
      RECT 146.09 95.7 147.41 95.9 ;
      RECT 146.09 97.62 147.41 97.82 ;
      RECT 146.09 99.1 147.41 99.3 ;
      RECT 146.09 101.02 147.41 101.22 ;
      RECT 146.09 102.5 147.41 102.7 ;
      RECT 146.09 104.42 147.41 104.62 ;
      RECT 146.09 105.9 147.41 106.1 ;
      RECT 146.09 107.82 147.41 108.02 ;
      RECT 146.09 109.3 147.41 109.5 ;
      RECT 146.09 111.22 147.41 111.42 ;
      RECT 146.09 112.7 147.41 112.9 ;
      RECT 146.09 114.62 147.41 114.82 ;
      RECT 146.09 116.1 147.41 116.3 ;
      RECT 146.09 118.02 147.41 118.22 ;
      RECT 146.09 119.5 147.41 119.7 ;
      RECT 146.09 121.42 147.41 121.62 ;
      RECT 146.09 122.9 147.41 123.1 ;
      RECT 146.09 124.82 147.41 125.02 ;
      RECT 146.09 126.3 147.41 126.5 ;
      RECT 146.09 128.22 147.41 128.42 ;
      RECT 146.09 129.7 147.41 129.9 ;
      RECT 146.09 131.62 147.41 131.82 ;
      RECT 146.09 133.1 147.41 133.3 ;
      RECT 146.09 135.02 147.41 135.22 ;
      RECT 146.09 136.5 147.41 136.7 ;
      RECT 146.09 138.42 147.41 138.62 ;
      RECT 146.09 139.9 147.41 140.1 ;
      RECT 146.09 141.82 147.41 142.02 ;
      RECT 146.09 143.3 147.41 143.5 ;
      RECT 146.09 145.22 147.41 145.42 ;
      RECT 146.09 146.7 147.41 146.9 ;
      RECT 146.09 148.62 147.41 148.82 ;
      RECT 146.09 150.1 147.41 150.3 ;
      RECT 146.09 152.02 147.41 152.22 ;
      RECT 146.09 153.5 147.41 153.7 ;
      RECT 146.09 155.42 147.41 155.62 ;
      RECT 146.09 156.9 147.41 157.1 ;
      RECT 146.09 158.82 147.41 159.02 ;
      RECT 146.09 160.3 147.41 160.5 ;
      RECT 146.09 162.22 147.41 162.42 ;
      RECT 146.09 163.7 147.41 163.9 ;
      RECT 146.09 165.62 147.41 165.82 ;
      RECT 146.09 167.1 147.41 167.3 ;
      RECT 146.09 169.02 147.41 169.22 ;
      RECT 146.09 170.5 147.41 170.7 ;
      RECT 146.09 172.42 147.41 172.62 ;
      RECT 146.09 173.9 147.41 174.1 ;
      RECT 146.09 175.82 147.41 176.02 ;
      RECT 146.09 177.3 147.41 177.5 ;
      RECT 146.09 179.22 147.41 179.42 ;
      RECT 146.09 180.7 147.41 180.9 ;
      RECT 146.09 182.62 147.41 182.82 ;
      RECT 146.09 184.1 147.41 184.3 ;
      RECT 146.09 186.02 147.41 186.22 ;
      RECT 146.09 187.5 147.41 187.7 ;
      RECT 146.09 189.42 147.41 189.62 ;
      RECT 146.09 190.9 147.41 191.1 ;
      RECT 146.09 192.82 147.41 193.02 ;
      RECT 146.09 194.3 147.41 194.5 ;
      RECT 146.09 196.22 147.41 196.42 ;
      RECT 146.09 197.7 147.41 197.9 ;
      RECT 146.09 199.62 147.41 199.82 ;
      RECT 146.09 201.1 147.41 201.3 ;
      RECT 146.09 203.02 147.41 203.22 ;
      RECT 146.09 204.5 147.41 204.7 ;
      RECT 146.09 206.42 147.41 206.62 ;
      RECT 146.09 207.9 147.41 208.1 ;
      RECT 146.09 209.82 147.41 210.02 ;
      RECT 146.09 211.3 147.41 211.5 ;
      RECT 146.09 213.22 147.41 213.42 ;
      RECT 146.09 214.7 147.41 214.9 ;
      RECT 146.09 216.62 147.41 216.82 ;
      RECT 146.09 218.1 147.41 218.3 ;
      RECT 146.09 220.02 147.41 220.22 ;
      RECT 146.09 221.5 147.41 221.7 ;
      RECT 146.09 223.42 147.41 223.62 ;
      RECT 146.09 224.9 147.41 225.1 ;
      RECT 146.09 226.82 147.41 227.02 ;
      RECT 146.09 228.3 147.41 228.5 ;
      RECT 146.09 230.22 147.41 230.42 ;
      RECT 146.09 231.7 147.41 231.9 ;
      RECT 146.09 233.62 147.41 233.82 ;
      RECT 146.09 235.1 147.41 235.3 ;
      RECT 146.09 237.02 147.41 237.22 ;
      RECT 146.09 238.5 147.41 238.7 ;
      RECT 146.09 240.42 147.41 240.62 ;
      RECT 146.09 241.9 147.41 242.1 ;
      RECT 146.09 243.82 147.41 244.02 ;
      RECT 146.09 245.3 147.41 245.5 ;
      RECT 146.09 247.22 147.41 247.42 ;
      RECT 146.09 248.7 147.41 248.9 ;
      RECT 146.09 250.62 147.41 250.82 ;
      RECT 146.09 252.1 147.41 252.3 ;
      RECT 146.09 254.02 147.41 254.22 ;
      RECT 146.09 255.5 147.41 255.7 ;
      RECT 146.09 257.42 147.41 257.62 ;
      RECT 146.09 258.9 147.41 259.1 ;
      RECT 146.09 260.82 147.41 261.02 ;
      RECT 146.09 262.3 147.41 262.5 ;
      RECT 146.09 264.22 147.41 264.42 ;
      RECT 146.09 265.7 147.41 265.9 ;
      RECT 146.09 267.62 147.41 267.82 ;
      RECT 146.09 269.1 147.41 269.3 ;
      RECT 146.09 271.02 147.41 271.22 ;
      RECT 146.09 272.5 147.41 272.7 ;
      RECT 146.09 274.42 147.41 274.62 ;
      RECT 146.09 275.9 147.41 276.1 ;
      RECT 146.09 277.82 147.41 278.02 ;
      RECT 146.09 279.3 147.41 279.5 ;
      RECT 146.09 281.22 147.41 281.42 ;
      RECT 146.09 282.7 147.41 282.9 ;
      RECT 146.09 284.62 147.41 284.82 ;
      RECT 146.09 286.1 147.41 286.3 ;
      RECT 146.09 288.02 147.41 288.22 ;
      RECT 146.09 289.5 147.41 289.7 ;
      RECT 146.09 291.42 147.41 291.62 ;
      RECT 146.09 292.9 147.41 293.1 ;
      RECT 146.09 294.82 147.41 295.02 ;
      RECT 146.09 296.3 147.41 296.5 ;
      RECT 146.09 298.22 147.41 298.42 ;
      RECT 146.09 299.7 147.41 299.9 ;
      RECT 146.09 301.62 147.41 301.82 ;
      RECT 146.09 303.1 147.41 303.3 ;
      RECT 146.09 305.02 147.41 305.22 ;
      RECT 146.09 306.5 147.41 306.7 ;
      RECT 146.09 308.42 147.41 308.62 ;
      RECT 146.09 309.9 147.41 310.1 ;
      RECT 146.09 311.82 147.41 312.02 ;
      RECT 146.09 313.3 147.41 313.5 ;
      RECT 146.09 315.22 147.41 315.42 ;
      RECT 146.09 316.7 147.41 316.9 ;
      RECT 146.09 318.62 147.41 318.82 ;
      RECT 146.09 320.1 147.41 320.3 ;
      RECT 146.09 322.02 147.41 322.22 ;
      RECT 146.09 323.5 147.41 323.7 ;
      RECT 146.09 325.42 147.41 325.62 ;
      RECT 146.09 326.9 147.41 327.1 ;
      RECT 146.09 328.82 147.41 329.02 ;
      RECT 146.09 330.3 147.41 330.5 ;
      RECT 146.09 332.22 147.41 332.42 ;
      RECT 146.09 333.7 147.41 333.9 ;
      RECT 146.09 335.62 147.41 335.82 ;
      RECT 146.09 337.1 147.41 337.3 ;
      RECT 146.09 339.02 147.41 339.22 ;
      RECT 146.09 340.5 147.41 340.7 ;
      RECT 146.09 342.42 147.41 342.62 ;
      RECT 146.09 343.9 147.41 344.1 ;
      RECT 146.09 345.82 147.41 346.02 ;
      RECT 146.09 347.3 147.41 347.5 ;
      RECT 146.09 349.22 147.41 349.42 ;
      RECT 146.09 350.7 147.41 350.9 ;
      RECT 146.09 352.62 147.41 352.82 ;
      RECT 146.09 354.1 147.41 354.3 ;
      RECT 146.09 356.02 147.41 356.22 ;
      RECT 146.09 357.5 147.41 357.7 ;
      RECT 146.09 359.42 147.41 359.62 ;
      RECT 146.09 360.9 147.41 361.1 ;
      RECT 146.09 362.82 147.41 363.02 ;
      RECT 146.09 364.3 147.41 364.5 ;
      RECT 146.09 366.22 147.41 366.42 ;
      RECT 146.09 367.7 147.41 367.9 ;
      RECT 146.09 369.62 147.41 369.82 ;
      RECT 146.09 371.1 147.41 371.3 ;
      RECT 146.09 373.02 147.41 373.22 ;
      RECT 146.09 374.5 147.41 374.7 ;
      RECT 146.09 376.42 147.41 376.62 ;
      RECT 146.09 377.9 147.41 378.1 ;
      RECT 146.09 379.82 147.41 380.02 ;
      RECT 146.09 381.3 147.41 381.5 ;
      RECT 146.09 383.22 147.41 383.42 ;
      RECT 146.09 384.7 147.41 384.9 ;
      RECT 146.09 386.62 147.41 386.82 ;
      RECT 146.09 388.1 147.41 388.3 ;
      RECT 146.09 390.02 147.41 390.22 ;
      RECT 146.09 391.5 147.41 391.7 ;
      RECT 146.09 393.42 147.41 393.62 ;
      RECT 146.09 394.9 147.41 395.1 ;
      RECT 146.09 396.82 147.41 397.02 ;
      RECT 146.09 398.3 147.41 398.5 ;
      RECT 146.09 400.22 147.41 400.42 ;
      RECT 146.09 401.7 147.41 401.9 ;
      RECT 146.09 403.62 147.41 403.82 ;
      RECT 146.09 405.1 147.41 405.3 ;
      RECT 146.09 407.02 147.41 407.22 ;
      RECT 146.09 408.5 147.41 408.7 ;
      RECT 146.09 410.42 147.41 410.62 ;
      RECT 146.09 411.9 147.41 412.1 ;
      RECT 146.09 413.82 147.41 414.02 ;
      RECT 146.09 415.3 147.41 415.5 ;
      RECT 146.09 417.22 147.41 417.42 ;
      RECT 146.09 418.7 147.41 418.9 ;
      RECT 146.09 420.62 147.41 420.82 ;
      RECT 146.09 422.1 147.41 422.3 ;
      RECT 146.09 424.02 147.41 424.22 ;
      RECT 146.09 425.5 147.41 425.7 ;
      RECT 146.09 427.42 147.41 427.62 ;
      RECT 146.09 428.9 147.41 429.1 ;
      RECT 146.09 430.82 147.41 431.02 ;
      RECT 146.09 432.3 147.41 432.5 ;
      RECT 146.09 434.22 147.41 434.42 ;
      RECT 146.09 435.7 147.41 435.9 ;
      RECT 146.09 437.62 147.41 437.82 ;
      RECT 146.09 439.1 147.41 439.3 ;
      RECT 146.09 441.02 147.41 441.22 ;
      RECT 146.09 442.5 147.41 442.7 ;
      RECT 146.09 444.42 147.41 444.62 ;
      RECT 146.09 445.9 147.41 446.1 ;
      RECT 146.09 447.82 147.41 448.02 ;
      RECT 146.09 449.3 147.41 449.5 ;
      RECT 146.09 451.22 147.41 451.42 ;
      RECT 146.09 452.7 147.41 452.9 ;
      RECT 146.09 454.62 147.41 454.82 ;
      RECT 146.09 456.1 147.41 456.3 ;
      RECT 146.09 458.02 147.41 458.22 ;
      RECT 146.09 459.5 147.41 459.7 ;
      RECT 146.09 461.42 147.41 461.62 ;
      RECT 146.09 462.9 147.41 463.1 ;
      RECT 146.09 464.82 147.41 465.02 ;
      RECT 146.09 466.3 147.41 466.5 ;
      RECT 146.09 468.22 147.41 468.42 ;
      RECT 146.09 469.7 147.41 469.9 ;
      RECT 146.09 471.62 147.41 471.82 ;
      RECT 146.09 473.1 147.41 473.3 ;
      RECT 146.09 475.02 147.41 475.22 ;
      RECT 146.09 476.5 147.41 476.7 ;
      RECT 146.09 478.42 147.41 478.62 ;
      RECT 146.09 479.9 147.41 480.1 ;
      RECT 146.09 481.82 147.41 482.02 ;
      RECT 146.09 483.3 147.41 483.5 ;
      RECT 146.09 485.22 147.41 485.42 ;
      RECT 146.09 486.7 147.41 486.9 ;
      RECT 146.09 488.62 147.41 488.82 ;
      RECT 146.09 490.1 147.41 490.3 ;
      RECT 146.09 492.02 147.41 492.22 ;
      RECT 146.09 493.5 147.41 493.7 ;
      RECT 146.09 495.42 147.41 495.62 ;
      RECT 146.09 496.9 147.41 497.1 ;
      RECT 146.09 498.82 147.41 499.02 ;
      RECT 146.09 500.3 147.41 500.5 ;
      RECT 146.09 502.22 147.41 502.42 ;
      RECT 146.09 503.7 147.41 503.9 ;
      RECT 146.09 505.62 147.41 505.82 ;
      RECT 146.09 510.34 147.41 510.94 ;
      RECT 145.13 29.53 147.39 29.73 ;
      RECT 144.26 29.93 146.99 30.13 ;
      RECT 145.06 52.16 146.54 52.76 ;
      RECT 145.65 62.18 145.93 62.78 ;
      RECT 145.01 6.24 145.61 6.84 ;
      RECT 144.17 510.34 145.49 510.94 ;
      RECT 144.21 10.23 145.45 10.83 ;
      RECT 143.12 52.16 144.6 52.76 ;
      RECT 143.81 16.74 144.35 17.34 ;
      RECT 142.52 29.64 144.01 29.84 ;
      RECT 143.73 62.18 144.01 62.78 ;
      RECT 142.62 6.24 143.57 6.84 ;
      RECT 142.25 510.34 143.57 510.94 ;
      RECT 141.22 52.16 142.7 52.76 ;
      RECT 141.62 6.24 142.22 6.84 ;
      RECT 141.99 29.37 142.22 30.28 ;
      RECT 141.81 62.18 142.09 62.78 ;
      RECT 138.41 510.34 141.65 510.94 ;
      RECT 135.81 70.42 141.63 70.62 ;
      RECT 135.81 71.9 141.63 72.1 ;
      RECT 135.81 73.82 141.63 74.02 ;
      RECT 135.81 75.3 141.63 75.5 ;
      RECT 135.81 77.22 141.63 77.42 ;
      RECT 135.81 78.7 141.63 78.9 ;
      RECT 135.81 80.62 141.63 80.82 ;
      RECT 135.81 82.1 141.63 82.3 ;
      RECT 135.81 84.02 141.63 84.22 ;
      RECT 135.81 85.5 141.63 85.7 ;
      RECT 135.81 87.42 141.63 87.62 ;
      RECT 135.81 88.9 141.63 89.1 ;
      RECT 135.81 90.82 141.63 91.02 ;
      RECT 135.81 92.3 141.63 92.5 ;
      RECT 135.81 94.22 141.63 94.42 ;
      RECT 135.81 95.7 141.63 95.9 ;
      RECT 135.81 97.62 141.63 97.82 ;
      RECT 135.81 99.1 141.63 99.3 ;
      RECT 135.81 101.02 141.63 101.22 ;
      RECT 135.81 102.5 141.63 102.7 ;
      RECT 135.81 104.42 141.63 104.62 ;
      RECT 135.81 105.9 141.63 106.1 ;
      RECT 135.81 107.82 141.63 108.02 ;
      RECT 135.81 109.3 141.63 109.5 ;
      RECT 135.81 111.22 141.63 111.42 ;
      RECT 135.81 112.7 141.63 112.9 ;
      RECT 135.81 114.62 141.63 114.82 ;
      RECT 135.81 116.1 141.63 116.3 ;
      RECT 135.81 118.02 141.63 118.22 ;
      RECT 135.81 119.5 141.63 119.7 ;
      RECT 135.81 121.42 141.63 121.62 ;
      RECT 135.81 122.9 141.63 123.1 ;
      RECT 135.81 124.82 141.63 125.02 ;
      RECT 135.81 126.3 141.63 126.5 ;
      RECT 135.81 128.22 141.63 128.42 ;
      RECT 135.81 129.7 141.63 129.9 ;
      RECT 135.81 131.62 141.63 131.82 ;
      RECT 135.81 133.1 141.63 133.3 ;
      RECT 135.81 135.02 141.63 135.22 ;
      RECT 135.81 136.5 141.63 136.7 ;
      RECT 135.81 138.42 141.63 138.62 ;
      RECT 135.81 139.9 141.63 140.1 ;
      RECT 135.81 141.82 141.63 142.02 ;
      RECT 135.81 143.3 141.63 143.5 ;
      RECT 135.81 145.22 141.63 145.42 ;
      RECT 135.81 146.7 141.63 146.9 ;
      RECT 135.81 148.62 141.63 148.82 ;
      RECT 135.81 150.1 141.63 150.3 ;
      RECT 135.81 152.02 141.63 152.22 ;
      RECT 135.81 153.5 141.63 153.7 ;
      RECT 135.81 155.42 141.63 155.62 ;
      RECT 135.81 156.9 141.63 157.1 ;
      RECT 135.81 158.82 141.63 159.02 ;
      RECT 135.81 160.3 141.63 160.5 ;
      RECT 135.81 162.22 141.63 162.42 ;
      RECT 135.81 163.7 141.63 163.9 ;
      RECT 135.81 165.62 141.63 165.82 ;
      RECT 135.81 167.1 141.63 167.3 ;
      RECT 135.81 169.02 141.63 169.22 ;
      RECT 135.81 170.5 141.63 170.7 ;
      RECT 135.81 172.42 141.63 172.62 ;
      RECT 135.81 173.9 141.63 174.1 ;
      RECT 135.81 175.82 141.63 176.02 ;
      RECT 135.81 177.3 141.63 177.5 ;
      RECT 135.81 179.22 141.63 179.42 ;
      RECT 135.81 180.7 141.63 180.9 ;
      RECT 135.81 182.62 141.63 182.82 ;
      RECT 135.81 184.1 141.63 184.3 ;
      RECT 135.81 186.02 141.63 186.22 ;
      RECT 135.81 187.5 141.63 187.7 ;
      RECT 135.81 189.42 141.63 189.62 ;
      RECT 135.81 190.9 141.63 191.1 ;
      RECT 135.81 192.82 141.63 193.02 ;
      RECT 135.81 194.3 141.63 194.5 ;
      RECT 135.81 196.22 141.63 196.42 ;
      RECT 135.81 197.7 141.63 197.9 ;
      RECT 135.81 199.62 141.63 199.82 ;
      RECT 135.81 201.1 141.63 201.3 ;
      RECT 135.81 203.02 141.63 203.22 ;
      RECT 135.81 204.5 141.63 204.7 ;
      RECT 135.81 206.42 141.63 206.62 ;
      RECT 135.81 207.9 141.63 208.1 ;
      RECT 135.81 209.82 141.63 210.02 ;
      RECT 135.81 211.3 141.63 211.5 ;
      RECT 135.81 213.22 141.63 213.42 ;
      RECT 135.81 214.7 141.63 214.9 ;
      RECT 135.81 216.62 141.63 216.82 ;
      RECT 135.81 218.1 141.63 218.3 ;
      RECT 135.81 220.02 141.63 220.22 ;
      RECT 135.81 221.5 141.63 221.7 ;
      RECT 135.81 223.42 141.63 223.62 ;
      RECT 135.81 224.9 141.63 225.1 ;
      RECT 135.81 226.82 141.63 227.02 ;
      RECT 135.81 228.3 141.63 228.5 ;
      RECT 135.81 230.22 141.63 230.42 ;
      RECT 135.81 231.7 141.63 231.9 ;
      RECT 135.81 233.62 141.63 233.82 ;
      RECT 135.81 235.1 141.63 235.3 ;
      RECT 135.81 237.02 141.63 237.22 ;
      RECT 135.81 238.5 141.63 238.7 ;
      RECT 135.81 240.42 141.63 240.62 ;
      RECT 135.81 241.9 141.63 242.1 ;
      RECT 135.81 243.82 141.63 244.02 ;
      RECT 135.81 245.3 141.63 245.5 ;
      RECT 135.81 247.22 141.63 247.42 ;
      RECT 135.81 248.7 141.63 248.9 ;
      RECT 135.81 250.62 141.63 250.82 ;
      RECT 135.81 252.1 141.63 252.3 ;
      RECT 135.81 254.02 141.63 254.22 ;
      RECT 135.81 255.5 141.63 255.7 ;
      RECT 135.81 257.42 141.63 257.62 ;
      RECT 135.81 258.9 141.63 259.1 ;
      RECT 135.81 260.82 141.63 261.02 ;
      RECT 135.81 262.3 141.63 262.5 ;
      RECT 135.81 264.22 141.63 264.42 ;
      RECT 135.81 265.7 141.63 265.9 ;
      RECT 135.81 267.62 141.63 267.82 ;
      RECT 135.81 269.1 141.63 269.3 ;
      RECT 135.81 271.02 141.63 271.22 ;
      RECT 135.81 272.5 141.63 272.7 ;
      RECT 135.81 274.42 141.63 274.62 ;
      RECT 135.81 275.9 141.63 276.1 ;
      RECT 135.81 277.82 141.63 278.02 ;
      RECT 135.81 279.3 141.63 279.5 ;
      RECT 135.81 281.22 141.63 281.42 ;
      RECT 135.81 282.7 141.63 282.9 ;
      RECT 135.81 284.62 141.63 284.82 ;
      RECT 135.81 286.1 141.63 286.3 ;
      RECT 135.81 288.02 141.63 288.22 ;
      RECT 135.81 289.5 141.63 289.7 ;
      RECT 135.81 291.42 141.63 291.62 ;
      RECT 135.81 292.9 141.63 293.1 ;
      RECT 135.81 294.82 141.63 295.02 ;
      RECT 135.81 296.3 141.63 296.5 ;
      RECT 135.81 298.22 141.63 298.42 ;
      RECT 135.81 299.7 141.63 299.9 ;
      RECT 135.81 301.62 141.63 301.82 ;
      RECT 135.81 303.1 141.63 303.3 ;
      RECT 135.81 305.02 141.63 305.22 ;
      RECT 135.81 306.5 141.63 306.7 ;
      RECT 135.81 308.42 141.63 308.62 ;
      RECT 135.81 309.9 141.63 310.1 ;
      RECT 135.81 311.82 141.63 312.02 ;
      RECT 135.81 313.3 141.63 313.5 ;
      RECT 135.81 315.22 141.63 315.42 ;
      RECT 135.81 316.7 141.63 316.9 ;
      RECT 135.81 318.62 141.63 318.82 ;
      RECT 135.81 320.1 141.63 320.3 ;
      RECT 135.81 322.02 141.63 322.22 ;
      RECT 135.81 323.5 141.63 323.7 ;
      RECT 135.81 325.42 141.63 325.62 ;
      RECT 135.81 326.9 141.63 327.1 ;
      RECT 135.81 328.82 141.63 329.02 ;
      RECT 135.81 330.3 141.63 330.5 ;
      RECT 135.81 332.22 141.63 332.42 ;
      RECT 135.81 333.7 141.63 333.9 ;
      RECT 135.81 335.62 141.63 335.82 ;
      RECT 135.81 337.1 141.63 337.3 ;
      RECT 135.81 339.02 141.63 339.22 ;
      RECT 135.81 340.5 141.63 340.7 ;
      RECT 135.81 342.42 141.63 342.62 ;
      RECT 135.81 343.9 141.63 344.1 ;
      RECT 135.81 345.82 141.63 346.02 ;
      RECT 135.81 347.3 141.63 347.5 ;
      RECT 135.81 349.22 141.63 349.42 ;
      RECT 135.81 350.7 141.63 350.9 ;
      RECT 135.81 352.62 141.63 352.82 ;
      RECT 135.81 354.1 141.63 354.3 ;
      RECT 135.81 356.02 141.63 356.22 ;
      RECT 135.81 357.5 141.63 357.7 ;
      RECT 135.81 359.42 141.63 359.62 ;
      RECT 135.81 360.9 141.63 361.1 ;
      RECT 135.81 362.82 141.63 363.02 ;
      RECT 135.81 364.3 141.63 364.5 ;
      RECT 135.81 366.22 141.63 366.42 ;
      RECT 135.81 367.7 141.63 367.9 ;
      RECT 135.81 369.62 141.63 369.82 ;
      RECT 135.81 371.1 141.63 371.3 ;
      RECT 135.81 373.02 141.63 373.22 ;
      RECT 135.81 374.5 141.63 374.7 ;
      RECT 135.81 376.42 141.63 376.62 ;
      RECT 135.81 377.9 141.63 378.1 ;
      RECT 135.81 379.82 141.63 380.02 ;
      RECT 135.81 381.3 141.63 381.5 ;
      RECT 135.81 383.22 141.63 383.42 ;
      RECT 135.81 384.7 141.63 384.9 ;
      RECT 135.81 386.62 141.63 386.82 ;
      RECT 135.81 388.1 141.63 388.3 ;
      RECT 135.81 390.02 141.63 390.22 ;
      RECT 135.81 391.5 141.63 391.7 ;
      RECT 135.81 393.42 141.63 393.62 ;
      RECT 135.81 394.9 141.63 395.1 ;
      RECT 135.81 396.82 141.63 397.02 ;
      RECT 135.81 398.3 141.63 398.5 ;
      RECT 135.81 400.22 141.63 400.42 ;
      RECT 135.81 401.7 141.63 401.9 ;
      RECT 135.81 403.62 141.63 403.82 ;
      RECT 135.81 405.1 141.63 405.3 ;
      RECT 135.81 407.02 141.63 407.22 ;
      RECT 135.81 408.5 141.63 408.7 ;
      RECT 135.81 410.42 141.63 410.62 ;
      RECT 135.81 411.9 141.63 412.1 ;
      RECT 135.81 413.82 141.63 414.02 ;
      RECT 135.81 415.3 141.63 415.5 ;
      RECT 135.81 417.22 141.63 417.42 ;
      RECT 135.81 418.7 141.63 418.9 ;
      RECT 135.81 420.62 141.63 420.82 ;
      RECT 135.81 422.1 141.63 422.3 ;
      RECT 135.81 424.02 141.63 424.22 ;
      RECT 135.81 425.5 141.63 425.7 ;
      RECT 135.81 427.42 141.63 427.62 ;
      RECT 135.81 428.9 141.63 429.1 ;
      RECT 135.81 430.82 141.63 431.02 ;
      RECT 135.81 432.3 141.63 432.5 ;
      RECT 135.81 434.22 141.63 434.42 ;
      RECT 135.81 435.7 141.63 435.9 ;
      RECT 135.81 437.62 141.63 437.82 ;
      RECT 135.81 439.1 141.63 439.3 ;
      RECT 135.81 441.02 141.63 441.22 ;
      RECT 135.81 442.5 141.63 442.7 ;
      RECT 135.81 444.42 141.63 444.62 ;
      RECT 135.81 445.9 141.63 446.1 ;
      RECT 135.81 447.82 141.63 448.02 ;
      RECT 135.81 449.3 141.63 449.5 ;
      RECT 135.81 451.22 141.63 451.42 ;
      RECT 135.81 452.7 141.63 452.9 ;
      RECT 135.81 454.62 141.63 454.82 ;
      RECT 135.81 456.1 141.63 456.3 ;
      RECT 135.81 458.02 141.63 458.22 ;
      RECT 135.81 459.5 141.63 459.7 ;
      RECT 135.81 461.42 141.63 461.62 ;
      RECT 135.81 462.9 141.63 463.1 ;
      RECT 135.81 464.82 141.63 465.02 ;
      RECT 135.81 466.3 141.63 466.5 ;
      RECT 135.81 468.22 141.63 468.42 ;
      RECT 135.81 469.7 141.63 469.9 ;
      RECT 135.81 471.62 141.63 471.82 ;
      RECT 135.81 473.1 141.63 473.3 ;
      RECT 135.81 475.02 141.63 475.22 ;
      RECT 135.81 476.5 141.63 476.7 ;
      RECT 135.81 478.42 141.63 478.62 ;
      RECT 135.81 479.9 141.63 480.1 ;
      RECT 135.81 481.82 141.63 482.02 ;
      RECT 135.81 483.3 141.63 483.5 ;
      RECT 135.81 485.22 141.63 485.42 ;
      RECT 135.81 486.7 141.63 486.9 ;
      RECT 135.81 488.62 141.63 488.82 ;
      RECT 135.81 490.1 141.63 490.3 ;
      RECT 135.81 492.02 141.63 492.22 ;
      RECT 135.81 493.5 141.63 493.7 ;
      RECT 135.81 495.42 141.63 495.62 ;
      RECT 135.81 496.9 141.63 497.1 ;
      RECT 135.81 498.82 141.63 499.02 ;
      RECT 135.81 500.3 141.63 500.5 ;
      RECT 135.81 502.22 141.63 502.42 ;
      RECT 135.81 503.7 141.63 503.9 ;
      RECT 138.83 6.24 140.83 6.84 ;
      RECT 88.21 24.03 140.41 24.43 ;
      RECT 88.21 57.62 140.41 58.02 ;
      RECT 87.61 42.78 139.91 43.78 ;
      RECT 138.41 12.32 139.43 12.52 ;
      RECT 137.09 30.6 139.17 30.8 ;
      RECT 137.09 51.44 139.17 51.64 ;
      RECT 138.01 12.82 139.09 13.02 ;
      RECT 138.41 37.58 138.72 38.38 ;
      RECT 138.01 16.13 138.21 16.73 ;
      RECT 138.01 62.01 138.21 62.79 ;
      RECT 136.79 13.78 137.81 13.98 ;
      RECT 137.41 37.58 137.81 38.38 ;
      RECT 135.01 510.34 137.81 510.94 ;
      RECT 135.43 6.24 137.39 6.84 ;
      RECT 135.01 13.78 136.03 13.98 ;
      RECT 133.65 30.6 135.73 30.8 ;
      RECT 133.65 51.44 135.73 51.64 ;
      RECT 124.81 35.33 135.21 35.53 ;
      RECT 133.73 12.82 134.81 13.02 ;
      RECT 134.61 16.13 134.81 16.73 ;
      RECT 134.61 62.01 134.81 62.79 ;
      RECT 133.39 12.32 134.41 12.52 ;
      RECT 130.81 34.53 134.41 34.73 ;
      RECT 134.1 37.58 134.41 38.38 ;
      RECT 131.61 70.42 134.41 70.62 ;
      RECT 131.61 71.9 134.41 72.1 ;
      RECT 131.61 73.82 134.41 74.02 ;
      RECT 131.61 75.3 134.41 75.5 ;
      RECT 131.61 77.22 134.41 77.42 ;
      RECT 131.61 78.7 134.41 78.9 ;
      RECT 131.61 80.62 134.41 80.82 ;
      RECT 131.61 82.1 134.41 82.3 ;
      RECT 131.61 84.02 134.41 84.22 ;
      RECT 131.61 85.5 134.41 85.7 ;
      RECT 131.61 87.42 134.41 87.62 ;
      RECT 131.61 88.9 134.41 89.1 ;
      RECT 131.61 90.82 134.41 91.02 ;
      RECT 131.61 92.3 134.41 92.5 ;
      RECT 131.61 94.22 134.41 94.42 ;
      RECT 131.61 95.7 134.41 95.9 ;
      RECT 131.61 97.62 134.41 97.82 ;
      RECT 131.61 99.1 134.41 99.3 ;
      RECT 131.61 101.02 134.41 101.22 ;
      RECT 131.61 102.5 134.41 102.7 ;
      RECT 131.61 104.42 134.41 104.62 ;
      RECT 131.61 105.9 134.41 106.1 ;
      RECT 131.61 107.82 134.41 108.02 ;
      RECT 131.61 109.3 134.41 109.5 ;
      RECT 131.61 111.22 134.41 111.42 ;
      RECT 131.61 112.7 134.41 112.9 ;
      RECT 131.61 114.62 134.41 114.82 ;
      RECT 131.61 116.1 134.41 116.3 ;
      RECT 131.61 118.02 134.41 118.22 ;
      RECT 131.61 119.5 134.41 119.7 ;
      RECT 131.61 121.42 134.41 121.62 ;
      RECT 131.61 122.9 134.41 123.1 ;
      RECT 131.61 124.82 134.41 125.02 ;
      RECT 131.61 126.3 134.41 126.5 ;
      RECT 131.61 128.22 134.41 128.42 ;
      RECT 131.61 129.7 134.41 129.9 ;
      RECT 131.61 131.62 134.41 131.82 ;
      RECT 131.61 133.1 134.41 133.3 ;
      RECT 131.61 135.02 134.41 135.22 ;
      RECT 131.61 136.5 134.41 136.7 ;
      RECT 131.61 138.42 134.41 138.62 ;
      RECT 131.61 139.9 134.41 140.1 ;
      RECT 131.61 141.82 134.41 142.02 ;
      RECT 131.61 143.3 134.41 143.5 ;
      RECT 131.61 145.22 134.41 145.42 ;
      RECT 131.61 146.7 134.41 146.9 ;
      RECT 131.61 148.62 134.41 148.82 ;
      RECT 131.61 150.1 134.41 150.3 ;
      RECT 131.61 152.02 134.41 152.22 ;
      RECT 131.61 153.5 134.41 153.7 ;
      RECT 131.61 155.42 134.41 155.62 ;
      RECT 131.61 156.9 134.41 157.1 ;
      RECT 131.61 158.82 134.41 159.02 ;
      RECT 131.61 160.3 134.41 160.5 ;
      RECT 131.61 162.22 134.41 162.42 ;
      RECT 131.61 163.7 134.41 163.9 ;
      RECT 131.61 165.62 134.41 165.82 ;
      RECT 131.61 167.1 134.41 167.3 ;
      RECT 131.61 169.02 134.41 169.22 ;
      RECT 131.61 170.5 134.41 170.7 ;
      RECT 131.61 172.42 134.41 172.62 ;
      RECT 131.61 173.9 134.41 174.1 ;
      RECT 131.61 175.82 134.41 176.02 ;
      RECT 131.61 177.3 134.41 177.5 ;
      RECT 131.61 179.22 134.41 179.42 ;
      RECT 131.61 180.7 134.41 180.9 ;
      RECT 131.61 182.62 134.41 182.82 ;
      RECT 131.61 184.1 134.41 184.3 ;
      RECT 131.61 186.02 134.41 186.22 ;
      RECT 131.61 187.5 134.41 187.7 ;
      RECT 131.61 189.42 134.41 189.62 ;
      RECT 131.61 190.9 134.41 191.1 ;
      RECT 131.61 192.82 134.41 193.02 ;
      RECT 131.61 194.3 134.41 194.5 ;
      RECT 131.61 196.22 134.41 196.42 ;
      RECT 131.61 197.7 134.41 197.9 ;
      RECT 131.61 199.62 134.41 199.82 ;
      RECT 131.61 201.1 134.41 201.3 ;
      RECT 131.61 203.02 134.41 203.22 ;
      RECT 131.61 204.5 134.41 204.7 ;
      RECT 131.61 206.42 134.41 206.62 ;
      RECT 131.61 207.9 134.41 208.1 ;
      RECT 131.61 209.82 134.41 210.02 ;
      RECT 131.61 211.3 134.41 211.5 ;
      RECT 131.61 213.22 134.41 213.42 ;
      RECT 131.61 214.7 134.41 214.9 ;
      RECT 131.61 216.62 134.41 216.82 ;
      RECT 131.61 218.1 134.41 218.3 ;
      RECT 131.61 220.02 134.41 220.22 ;
      RECT 131.61 221.5 134.41 221.7 ;
      RECT 131.61 223.42 134.41 223.62 ;
      RECT 131.61 224.9 134.41 225.1 ;
      RECT 131.61 226.82 134.41 227.02 ;
      RECT 131.61 228.3 134.41 228.5 ;
      RECT 131.61 230.22 134.41 230.42 ;
      RECT 131.61 231.7 134.41 231.9 ;
      RECT 131.61 233.62 134.41 233.82 ;
      RECT 131.61 235.1 134.41 235.3 ;
      RECT 131.61 237.02 134.41 237.22 ;
      RECT 131.61 238.5 134.41 238.7 ;
      RECT 131.61 240.42 134.41 240.62 ;
      RECT 131.61 241.9 134.41 242.1 ;
      RECT 131.61 243.82 134.41 244.02 ;
      RECT 131.61 245.3 134.41 245.5 ;
      RECT 131.61 247.22 134.41 247.42 ;
      RECT 131.61 248.7 134.41 248.9 ;
      RECT 131.61 250.62 134.41 250.82 ;
      RECT 131.61 252.1 134.41 252.3 ;
      RECT 131.61 254.02 134.41 254.22 ;
      RECT 131.61 255.5 134.41 255.7 ;
      RECT 131.61 257.42 134.41 257.62 ;
      RECT 131.61 258.9 134.41 259.1 ;
      RECT 131.61 260.82 134.41 261.02 ;
      RECT 131.61 262.3 134.41 262.5 ;
      RECT 131.61 264.22 134.41 264.42 ;
      RECT 131.61 265.7 134.41 265.9 ;
      RECT 131.61 267.62 134.41 267.82 ;
      RECT 131.61 269.1 134.41 269.3 ;
      RECT 131.61 271.02 134.41 271.22 ;
      RECT 131.61 272.5 134.41 272.7 ;
      RECT 131.61 274.42 134.41 274.62 ;
      RECT 131.61 275.9 134.41 276.1 ;
      RECT 131.61 277.82 134.41 278.02 ;
      RECT 131.61 279.3 134.41 279.5 ;
      RECT 131.61 281.22 134.41 281.42 ;
      RECT 131.61 282.7 134.41 282.9 ;
      RECT 131.61 284.62 134.41 284.82 ;
      RECT 131.61 286.1 134.41 286.3 ;
      RECT 131.61 288.02 134.41 288.22 ;
      RECT 131.61 289.5 134.41 289.7 ;
      RECT 131.61 291.42 134.41 291.62 ;
      RECT 131.61 292.9 134.41 293.1 ;
      RECT 131.61 294.82 134.41 295.02 ;
      RECT 131.61 296.3 134.41 296.5 ;
      RECT 131.61 298.22 134.41 298.42 ;
      RECT 131.61 299.7 134.41 299.9 ;
      RECT 131.61 301.62 134.41 301.82 ;
      RECT 131.61 303.1 134.41 303.3 ;
      RECT 131.61 305.02 134.41 305.22 ;
      RECT 131.61 306.5 134.41 306.7 ;
      RECT 131.61 308.42 134.41 308.62 ;
      RECT 131.61 309.9 134.41 310.1 ;
      RECT 131.61 311.82 134.41 312.02 ;
      RECT 131.61 313.3 134.41 313.5 ;
      RECT 131.61 315.22 134.41 315.42 ;
      RECT 131.61 316.7 134.41 316.9 ;
      RECT 131.61 318.62 134.41 318.82 ;
      RECT 131.61 320.1 134.41 320.3 ;
      RECT 131.61 322.02 134.41 322.22 ;
      RECT 131.61 323.5 134.41 323.7 ;
      RECT 131.61 325.42 134.41 325.62 ;
      RECT 131.61 326.9 134.41 327.1 ;
      RECT 131.61 328.82 134.41 329.02 ;
      RECT 131.61 330.3 134.41 330.5 ;
      RECT 131.61 332.22 134.41 332.42 ;
      RECT 131.61 333.7 134.41 333.9 ;
      RECT 131.61 335.62 134.41 335.82 ;
      RECT 131.61 337.1 134.41 337.3 ;
      RECT 131.61 339.02 134.41 339.22 ;
      RECT 131.61 340.5 134.41 340.7 ;
      RECT 131.61 342.42 134.41 342.62 ;
      RECT 131.61 343.9 134.41 344.1 ;
      RECT 131.61 345.82 134.41 346.02 ;
      RECT 131.61 347.3 134.41 347.5 ;
      RECT 131.61 349.22 134.41 349.42 ;
      RECT 131.61 350.7 134.41 350.9 ;
      RECT 131.61 352.62 134.41 352.82 ;
      RECT 131.61 354.1 134.41 354.3 ;
      RECT 131.61 356.02 134.41 356.22 ;
      RECT 131.61 357.5 134.41 357.7 ;
      RECT 131.61 359.42 134.41 359.62 ;
      RECT 131.61 360.9 134.41 361.1 ;
      RECT 131.61 362.82 134.41 363.02 ;
      RECT 131.61 364.3 134.41 364.5 ;
      RECT 131.61 366.22 134.41 366.42 ;
      RECT 131.61 367.7 134.41 367.9 ;
      RECT 131.61 369.62 134.41 369.82 ;
      RECT 131.61 371.1 134.41 371.3 ;
      RECT 131.61 373.02 134.41 373.22 ;
      RECT 131.61 374.5 134.41 374.7 ;
      RECT 131.61 376.42 134.41 376.62 ;
      RECT 131.61 377.9 134.41 378.1 ;
      RECT 131.61 379.82 134.41 380.02 ;
      RECT 131.61 381.3 134.41 381.5 ;
      RECT 131.61 383.22 134.41 383.42 ;
      RECT 131.61 384.7 134.41 384.9 ;
      RECT 131.61 386.62 134.41 386.82 ;
      RECT 131.61 388.1 134.41 388.3 ;
      RECT 131.61 390.02 134.41 390.22 ;
      RECT 131.61 391.5 134.41 391.7 ;
      RECT 131.61 393.42 134.41 393.62 ;
      RECT 131.61 394.9 134.41 395.1 ;
      RECT 131.61 396.82 134.41 397.02 ;
      RECT 131.61 398.3 134.41 398.5 ;
      RECT 131.61 400.22 134.41 400.42 ;
      RECT 131.61 401.7 134.41 401.9 ;
      RECT 131.61 403.62 134.41 403.82 ;
      RECT 131.61 405.1 134.41 405.3 ;
      RECT 131.61 407.02 134.41 407.22 ;
      RECT 131.61 408.5 134.41 408.7 ;
      RECT 131.61 410.42 134.41 410.62 ;
      RECT 131.61 411.9 134.41 412.1 ;
      RECT 131.61 413.82 134.41 414.02 ;
      RECT 131.61 415.3 134.41 415.5 ;
      RECT 131.61 417.22 134.41 417.42 ;
      RECT 131.61 418.7 134.41 418.9 ;
      RECT 131.61 420.62 134.41 420.82 ;
      RECT 131.61 422.1 134.41 422.3 ;
      RECT 131.61 424.02 134.41 424.22 ;
      RECT 131.61 425.5 134.41 425.7 ;
      RECT 131.61 427.42 134.41 427.62 ;
      RECT 131.61 428.9 134.41 429.1 ;
      RECT 131.61 430.82 134.41 431.02 ;
      RECT 131.61 432.3 134.41 432.5 ;
      RECT 131.61 434.22 134.41 434.42 ;
      RECT 131.61 435.7 134.41 435.9 ;
      RECT 131.61 437.62 134.41 437.82 ;
      RECT 131.61 439.1 134.41 439.3 ;
      RECT 131.61 441.02 134.41 441.22 ;
      RECT 131.61 442.5 134.41 442.7 ;
      RECT 131.61 444.42 134.41 444.62 ;
      RECT 131.61 445.9 134.41 446.1 ;
      RECT 131.61 447.82 134.41 448.02 ;
      RECT 131.61 449.3 134.41 449.5 ;
      RECT 131.61 451.22 134.41 451.42 ;
      RECT 131.61 452.7 134.41 452.9 ;
      RECT 131.61 454.62 134.41 454.82 ;
      RECT 131.61 456.1 134.41 456.3 ;
      RECT 131.61 458.02 134.41 458.22 ;
      RECT 131.61 459.5 134.41 459.7 ;
      RECT 131.61 461.42 134.41 461.62 ;
      RECT 131.61 462.9 134.41 463.1 ;
      RECT 131.61 464.82 134.41 465.02 ;
      RECT 131.61 466.3 134.41 466.5 ;
      RECT 131.61 468.22 134.41 468.42 ;
      RECT 131.61 469.7 134.41 469.9 ;
      RECT 131.61 471.62 134.41 471.82 ;
      RECT 131.61 473.1 134.41 473.3 ;
      RECT 131.61 475.02 134.41 475.22 ;
      RECT 131.61 476.5 134.41 476.7 ;
      RECT 131.61 478.42 134.41 478.62 ;
      RECT 131.61 479.9 134.41 480.1 ;
      RECT 131.61 481.82 134.41 482.02 ;
      RECT 131.61 483.3 134.41 483.5 ;
      RECT 131.61 485.22 134.41 485.42 ;
      RECT 131.61 486.7 134.41 486.9 ;
      RECT 131.61 488.62 134.41 488.82 ;
      RECT 131.61 490.1 134.41 490.3 ;
      RECT 131.61 492.02 134.41 492.22 ;
      RECT 131.61 493.5 134.41 493.7 ;
      RECT 131.61 495.42 134.41 495.62 ;
      RECT 131.61 496.9 134.41 497.1 ;
      RECT 131.61 498.82 134.41 499.02 ;
      RECT 131.61 500.3 134.41 500.5 ;
      RECT 131.61 502.22 134.41 502.42 ;
      RECT 131.61 503.7 134.41 503.9 ;
      RECT 131.61 510.34 134.41 510.94 ;
      RECT 111.06 508.84 134.01 509.04 ;
      RECT 132.03 6.24 133.99 6.84 ;
      RECT 126.9 32.48 133.9 32.68 ;
      RECT 133.7 37.58 133.9 38.38 ;
      RECT 124.73 506.34 133.61 506.54 ;
      RECT 131.61 12.32 132.63 12.52 ;
      RECT 130.29 30.6 132.37 30.8 ;
      RECT 130.29 51.44 132.37 51.64 ;
      RECT 125.31 34.93 132.32 35.13 ;
      RECT 132.12 37.58 132.32 38.38 ;
      RECT 131.21 12.82 132.29 13.02 ;
      RECT 131.61 37.58 131.92 38.38 ;
      RECT 131.21 16.13 131.41 16.73 ;
      RECT 131.21 62.01 131.41 62.79 ;
      RECT 129.99 13.78 131.01 13.98 ;
      RECT 128.21 69.46 131.01 69.66 ;
      RECT 128.21 72.86 131.01 73.06 ;
      RECT 128.21 76.26 131.01 76.46 ;
      RECT 128.21 79.66 131.01 79.86 ;
      RECT 128.21 83.06 131.01 83.26 ;
      RECT 128.21 86.46 131.01 86.66 ;
      RECT 128.21 89.86 131.01 90.06 ;
      RECT 128.21 93.26 131.01 93.46 ;
      RECT 128.21 96.66 131.01 96.86 ;
      RECT 128.21 100.06 131.01 100.26 ;
      RECT 128.21 103.46 131.01 103.66 ;
      RECT 128.21 106.86 131.01 107.06 ;
      RECT 128.21 110.26 131.01 110.46 ;
      RECT 128.21 113.66 131.01 113.86 ;
      RECT 128.21 117.06 131.01 117.26 ;
      RECT 128.21 120.46 131.01 120.66 ;
      RECT 128.21 123.86 131.01 124.06 ;
      RECT 128.21 127.26 131.01 127.46 ;
      RECT 128.21 130.66 131.01 130.86 ;
      RECT 128.21 134.06 131.01 134.26 ;
      RECT 128.21 137.46 131.01 137.66 ;
      RECT 128.21 140.86 131.01 141.06 ;
      RECT 128.21 144.26 131.01 144.46 ;
      RECT 128.21 147.66 131.01 147.86 ;
      RECT 128.21 151.06 131.01 151.26 ;
      RECT 128.21 154.46 131.01 154.66 ;
      RECT 128.21 157.86 131.01 158.06 ;
      RECT 128.21 161.26 131.01 161.46 ;
      RECT 128.21 164.66 131.01 164.86 ;
      RECT 128.21 168.06 131.01 168.26 ;
      RECT 128.21 171.46 131.01 171.66 ;
      RECT 128.21 174.86 131.01 175.06 ;
      RECT 128.21 178.26 131.01 178.46 ;
      RECT 128.21 181.66 131.01 181.86 ;
      RECT 128.21 185.06 131.01 185.26 ;
      RECT 128.21 188.46 131.01 188.66 ;
      RECT 128.21 191.86 131.01 192.06 ;
      RECT 128.21 195.26 131.01 195.46 ;
      RECT 128.21 198.66 131.01 198.86 ;
      RECT 128.21 202.06 131.01 202.26 ;
      RECT 128.21 205.46 131.01 205.66 ;
      RECT 128.21 208.86 131.01 209.06 ;
      RECT 128.21 212.26 131.01 212.46 ;
      RECT 128.21 215.66 131.01 215.86 ;
      RECT 128.21 219.06 131.01 219.26 ;
      RECT 128.21 222.46 131.01 222.66 ;
      RECT 128.21 225.86 131.01 226.06 ;
      RECT 128.21 229.26 131.01 229.46 ;
      RECT 128.21 232.66 131.01 232.86 ;
      RECT 128.21 236.06 131.01 236.26 ;
      RECT 128.21 239.46 131.01 239.66 ;
      RECT 128.21 242.86 131.01 243.06 ;
      RECT 128.21 246.26 131.01 246.46 ;
      RECT 128.21 249.66 131.01 249.86 ;
      RECT 128.21 253.06 131.01 253.26 ;
      RECT 128.21 256.46 131.01 256.66 ;
      RECT 128.21 259.86 131.01 260.06 ;
      RECT 128.21 263.26 131.01 263.46 ;
      RECT 128.21 266.66 131.01 266.86 ;
      RECT 128.21 270.06 131.01 270.26 ;
      RECT 128.21 273.46 131.01 273.66 ;
      RECT 128.21 276.86 131.01 277.06 ;
      RECT 128.21 280.26 131.01 280.46 ;
      RECT 128.21 283.66 131.01 283.86 ;
      RECT 128.21 287.06 131.01 287.26 ;
      RECT 128.21 290.46 131.01 290.66 ;
      RECT 128.21 293.86 131.01 294.06 ;
      RECT 128.21 297.26 131.01 297.46 ;
      RECT 128.21 300.66 131.01 300.86 ;
      RECT 128.21 304.06 131.01 304.26 ;
      RECT 128.21 307.46 131.01 307.66 ;
      RECT 128.21 310.86 131.01 311.06 ;
      RECT 128.21 314.26 131.01 314.46 ;
      RECT 128.21 317.66 131.01 317.86 ;
      RECT 128.21 321.06 131.01 321.26 ;
      RECT 128.21 324.46 131.01 324.66 ;
      RECT 128.21 327.86 131.01 328.06 ;
      RECT 128.21 331.26 131.01 331.46 ;
      RECT 128.21 334.66 131.01 334.86 ;
      RECT 128.21 338.06 131.01 338.26 ;
      RECT 128.21 341.46 131.01 341.66 ;
      RECT 128.21 344.86 131.01 345.06 ;
      RECT 128.21 348.26 131.01 348.46 ;
      RECT 128.21 351.66 131.01 351.86 ;
      RECT 128.21 355.06 131.01 355.26 ;
      RECT 128.21 358.46 131.01 358.66 ;
      RECT 128.21 361.86 131.01 362.06 ;
      RECT 128.21 365.26 131.01 365.46 ;
      RECT 128.21 368.66 131.01 368.86 ;
      RECT 128.21 372.06 131.01 372.26 ;
      RECT 128.21 375.46 131.01 375.66 ;
      RECT 128.21 378.86 131.01 379.06 ;
      RECT 128.21 382.26 131.01 382.46 ;
      RECT 128.21 385.66 131.01 385.86 ;
      RECT 128.21 389.06 131.01 389.26 ;
      RECT 128.21 392.46 131.01 392.66 ;
      RECT 128.21 395.86 131.01 396.06 ;
      RECT 128.21 399.26 131.01 399.46 ;
      RECT 128.21 402.66 131.01 402.86 ;
      RECT 128.21 406.06 131.01 406.26 ;
      RECT 128.21 409.46 131.01 409.66 ;
      RECT 128.21 412.86 131.01 413.06 ;
      RECT 128.21 416.26 131.01 416.46 ;
      RECT 128.21 419.66 131.01 419.86 ;
      RECT 128.21 423.06 131.01 423.26 ;
      RECT 128.21 426.46 131.01 426.66 ;
      RECT 128.21 429.86 131.01 430.06 ;
      RECT 128.21 433.26 131.01 433.46 ;
      RECT 128.21 436.66 131.01 436.86 ;
      RECT 128.21 440.06 131.01 440.26 ;
      RECT 128.21 443.46 131.01 443.66 ;
      RECT 128.21 446.86 131.01 447.06 ;
      RECT 128.21 450.26 131.01 450.46 ;
      RECT 128.21 453.66 131.01 453.86 ;
      RECT 128.21 457.06 131.01 457.26 ;
      RECT 128.21 460.46 131.01 460.66 ;
      RECT 128.21 463.86 131.01 464.06 ;
      RECT 128.21 467.26 131.01 467.46 ;
      RECT 128.21 470.66 131.01 470.86 ;
      RECT 128.21 474.06 131.01 474.26 ;
      RECT 128.21 477.46 131.01 477.66 ;
      RECT 128.21 480.86 131.01 481.06 ;
      RECT 128.21 484.26 131.01 484.46 ;
      RECT 128.21 487.66 131.01 487.86 ;
      RECT 128.21 491.06 131.01 491.26 ;
      RECT 128.21 494.46 131.01 494.66 ;
      RECT 128.21 497.86 131.01 498.06 ;
      RECT 128.21 501.26 131.01 501.46 ;
      RECT 128.21 504.66 131.01 504.86 ;
      RECT 128.21 510.34 131.01 510.94 ;
      RECT 128.63 6.24 130.59 6.84 ;
      RECT 128.21 34.53 130.4 34.73 ;
      RECT 123.22 70.36 129.66 70.56 ;
      RECT 123.22 71.96 129.66 72.16 ;
      RECT 123.22 73.76 129.66 73.96 ;
      RECT 123.22 75.36 129.66 75.56 ;
      RECT 123.22 77.16 129.66 77.36 ;
      RECT 123.22 78.76 129.66 78.96 ;
      RECT 123.22 80.56 129.66 80.76 ;
      RECT 123.22 82.16 129.66 82.36 ;
      RECT 123.22 83.96 129.66 84.16 ;
      RECT 123.22 85.56 129.66 85.76 ;
      RECT 123.22 87.36 129.66 87.56 ;
      RECT 123.22 88.96 129.66 89.16 ;
      RECT 123.22 90.76 129.66 90.96 ;
      RECT 123.22 92.36 129.66 92.56 ;
      RECT 123.22 94.16 129.66 94.36 ;
      RECT 123.22 95.76 129.66 95.96 ;
      RECT 123.22 97.56 129.66 97.76 ;
      RECT 123.22 99.16 129.66 99.36 ;
      RECT 123.22 100.96 129.66 101.16 ;
      RECT 123.22 102.56 129.66 102.76 ;
      RECT 123.22 104.36 129.66 104.56 ;
      RECT 123.22 105.96 129.66 106.16 ;
      RECT 123.22 107.76 129.66 107.96 ;
      RECT 123.22 109.36 129.66 109.56 ;
      RECT 123.22 111.16 129.66 111.36 ;
      RECT 123.22 112.76 129.66 112.96 ;
      RECT 123.22 114.56 129.66 114.76 ;
      RECT 123.22 116.16 129.66 116.36 ;
      RECT 123.22 117.96 129.66 118.16 ;
      RECT 123.22 119.56 129.66 119.76 ;
      RECT 123.22 121.36 129.66 121.56 ;
      RECT 123.22 122.96 129.66 123.16 ;
      RECT 123.22 124.76 129.66 124.96 ;
      RECT 123.22 126.36 129.66 126.56 ;
      RECT 123.22 128.16 129.66 128.36 ;
      RECT 123.22 129.76 129.66 129.96 ;
      RECT 123.22 131.56 129.66 131.76 ;
      RECT 123.22 133.16 129.66 133.36 ;
      RECT 123.22 134.96 129.66 135.16 ;
      RECT 123.22 136.56 129.66 136.76 ;
      RECT 123.22 138.36 129.66 138.56 ;
      RECT 123.22 139.96 129.66 140.16 ;
      RECT 123.22 141.76 129.66 141.96 ;
      RECT 123.22 143.36 129.66 143.56 ;
      RECT 123.22 145.16 129.66 145.36 ;
      RECT 123.22 146.76 129.66 146.96 ;
      RECT 123.22 148.56 129.66 148.76 ;
      RECT 123.22 150.16 129.66 150.36 ;
      RECT 123.22 151.96 129.66 152.16 ;
      RECT 123.22 153.56 129.66 153.76 ;
      RECT 123.22 155.36 129.66 155.56 ;
      RECT 123.22 156.96 129.66 157.16 ;
      RECT 123.22 158.76 129.66 158.96 ;
      RECT 123.22 160.36 129.66 160.56 ;
      RECT 123.22 162.16 129.66 162.36 ;
      RECT 123.22 163.76 129.66 163.96 ;
      RECT 123.22 165.56 129.66 165.76 ;
      RECT 123.22 167.16 129.66 167.36 ;
      RECT 123.22 168.96 129.66 169.16 ;
      RECT 123.22 170.56 129.66 170.76 ;
      RECT 123.22 172.36 129.66 172.56 ;
      RECT 123.22 173.96 129.66 174.16 ;
      RECT 123.22 175.76 129.66 175.96 ;
      RECT 123.22 177.36 129.66 177.56 ;
      RECT 123.22 179.16 129.66 179.36 ;
      RECT 123.22 180.76 129.66 180.96 ;
      RECT 123.22 182.56 129.66 182.76 ;
      RECT 123.22 184.16 129.66 184.36 ;
      RECT 123.22 185.96 129.66 186.16 ;
      RECT 123.22 187.56 129.66 187.76 ;
      RECT 123.22 189.36 129.66 189.56 ;
      RECT 123.22 190.96 129.66 191.16 ;
      RECT 123.22 192.76 129.66 192.96 ;
      RECT 123.22 194.36 129.66 194.56 ;
      RECT 123.22 196.16 129.66 196.36 ;
      RECT 123.22 197.76 129.66 197.96 ;
      RECT 123.22 199.56 129.66 199.76 ;
      RECT 123.22 201.16 129.66 201.36 ;
      RECT 123.22 202.96 129.66 203.16 ;
      RECT 123.22 204.56 129.66 204.76 ;
      RECT 123.22 206.36 129.66 206.56 ;
      RECT 123.22 207.96 129.66 208.16 ;
      RECT 123.22 209.76 129.66 209.96 ;
      RECT 123.22 211.36 129.66 211.56 ;
      RECT 123.22 213.16 129.66 213.36 ;
      RECT 123.22 214.76 129.66 214.96 ;
      RECT 123.22 216.56 129.66 216.76 ;
      RECT 123.22 218.16 129.66 218.36 ;
      RECT 123.22 219.96 129.66 220.16 ;
      RECT 123.22 221.56 129.66 221.76 ;
      RECT 123.22 223.36 129.66 223.56 ;
      RECT 123.22 224.96 129.66 225.16 ;
      RECT 123.22 226.76 129.66 226.96 ;
      RECT 123.22 228.36 129.66 228.56 ;
      RECT 123.22 230.16 129.66 230.36 ;
      RECT 123.22 231.76 129.66 231.96 ;
      RECT 123.22 233.56 129.66 233.76 ;
      RECT 123.22 235.16 129.66 235.36 ;
      RECT 123.22 236.96 129.66 237.16 ;
      RECT 123.22 238.56 129.66 238.76 ;
      RECT 123.22 240.36 129.66 240.56 ;
      RECT 123.22 241.96 129.66 242.16 ;
      RECT 123.22 243.76 129.66 243.96 ;
      RECT 123.22 245.36 129.66 245.56 ;
      RECT 123.22 247.16 129.66 247.36 ;
      RECT 123.22 248.76 129.66 248.96 ;
      RECT 123.22 250.56 129.66 250.76 ;
      RECT 123.22 252.16 129.66 252.36 ;
      RECT 123.22 253.96 129.66 254.16 ;
      RECT 123.22 255.56 129.66 255.76 ;
      RECT 123.22 257.36 129.66 257.56 ;
      RECT 123.22 258.96 129.66 259.16 ;
      RECT 123.22 260.76 129.66 260.96 ;
      RECT 123.22 262.36 129.66 262.56 ;
      RECT 123.22 264.16 129.66 264.36 ;
      RECT 123.22 265.76 129.66 265.96 ;
      RECT 123.22 267.56 129.66 267.76 ;
      RECT 123.22 269.16 129.66 269.36 ;
      RECT 123.22 270.96 129.66 271.16 ;
      RECT 123.22 272.56 129.66 272.76 ;
      RECT 123.22 274.36 129.66 274.56 ;
      RECT 123.22 275.96 129.66 276.16 ;
      RECT 123.22 277.76 129.66 277.96 ;
      RECT 123.22 279.36 129.66 279.56 ;
      RECT 123.22 281.16 129.66 281.36 ;
      RECT 123.22 282.76 129.66 282.96 ;
      RECT 123.22 284.56 129.66 284.76 ;
      RECT 123.22 286.16 129.66 286.36 ;
      RECT 123.22 287.96 129.66 288.16 ;
      RECT 123.22 289.56 129.66 289.76 ;
      RECT 123.22 291.36 129.66 291.56 ;
      RECT 123.22 292.96 129.66 293.16 ;
      RECT 123.22 294.76 129.66 294.96 ;
      RECT 123.22 296.36 129.66 296.56 ;
      RECT 123.22 298.16 129.66 298.36 ;
      RECT 123.22 299.76 129.66 299.96 ;
      RECT 123.22 301.56 129.66 301.76 ;
      RECT 123.22 303.16 129.66 303.36 ;
      RECT 123.22 304.96 129.66 305.16 ;
      RECT 123.22 306.56 129.66 306.76 ;
      RECT 123.22 308.36 129.66 308.56 ;
      RECT 123.22 309.96 129.66 310.16 ;
      RECT 123.22 311.76 129.66 311.96 ;
      RECT 123.22 313.36 129.66 313.56 ;
      RECT 123.22 315.16 129.66 315.36 ;
      RECT 123.22 316.76 129.66 316.96 ;
      RECT 123.22 318.56 129.66 318.76 ;
      RECT 123.22 320.16 129.66 320.36 ;
      RECT 123.22 321.96 129.66 322.16 ;
      RECT 123.22 323.56 129.66 323.76 ;
      RECT 123.22 325.36 129.66 325.56 ;
      RECT 123.22 326.96 129.66 327.16 ;
      RECT 123.22 328.76 129.66 328.96 ;
      RECT 123.22 330.36 129.66 330.56 ;
      RECT 123.22 332.16 129.66 332.36 ;
      RECT 123.22 333.76 129.66 333.96 ;
      RECT 123.22 335.56 129.66 335.76 ;
      RECT 123.22 337.16 129.66 337.36 ;
      RECT 123.22 338.96 129.66 339.16 ;
      RECT 123.22 340.56 129.66 340.76 ;
      RECT 123.22 342.36 129.66 342.56 ;
      RECT 123.22 343.96 129.66 344.16 ;
      RECT 123.22 345.76 129.66 345.96 ;
      RECT 123.22 347.36 129.66 347.56 ;
      RECT 123.22 349.16 129.66 349.36 ;
      RECT 123.22 350.76 129.66 350.96 ;
      RECT 123.22 352.56 129.66 352.76 ;
      RECT 123.22 354.16 129.66 354.36 ;
      RECT 123.22 355.96 129.66 356.16 ;
      RECT 123.22 357.56 129.66 357.76 ;
      RECT 123.22 359.36 129.66 359.56 ;
      RECT 123.22 360.96 129.66 361.16 ;
      RECT 123.22 362.76 129.66 362.96 ;
      RECT 123.22 364.36 129.66 364.56 ;
      RECT 123.22 366.16 129.66 366.36 ;
      RECT 123.22 367.76 129.66 367.96 ;
      RECT 123.22 369.56 129.66 369.76 ;
      RECT 123.22 371.16 129.66 371.36 ;
      RECT 123.22 372.96 129.66 373.16 ;
      RECT 123.22 374.56 129.66 374.76 ;
      RECT 123.22 376.36 129.66 376.56 ;
      RECT 123.22 377.96 129.66 378.16 ;
      RECT 123.22 379.76 129.66 379.96 ;
      RECT 123.22 381.36 129.66 381.56 ;
      RECT 123.22 383.16 129.66 383.36 ;
      RECT 123.22 384.76 129.66 384.96 ;
      RECT 123.22 386.56 129.66 386.76 ;
      RECT 123.22 388.16 129.66 388.36 ;
      RECT 123.22 389.96 129.66 390.16 ;
      RECT 123.22 391.56 129.66 391.76 ;
      RECT 123.22 393.36 129.66 393.56 ;
      RECT 123.22 394.96 129.66 395.16 ;
      RECT 123.22 396.76 129.66 396.96 ;
      RECT 123.22 398.36 129.66 398.56 ;
      RECT 123.22 400.16 129.66 400.36 ;
      RECT 123.22 401.76 129.66 401.96 ;
      RECT 123.22 403.56 129.66 403.76 ;
      RECT 123.22 405.16 129.66 405.36 ;
      RECT 123.22 406.96 129.66 407.16 ;
      RECT 123.22 408.56 129.66 408.76 ;
      RECT 123.22 410.36 129.66 410.56 ;
      RECT 123.22 411.96 129.66 412.16 ;
      RECT 123.22 413.76 129.66 413.96 ;
      RECT 123.22 415.36 129.66 415.56 ;
      RECT 123.22 417.16 129.66 417.36 ;
      RECT 123.22 418.76 129.66 418.96 ;
      RECT 123.22 420.56 129.66 420.76 ;
      RECT 123.22 422.16 129.66 422.36 ;
      RECT 123.22 423.96 129.66 424.16 ;
      RECT 123.22 425.56 129.66 425.76 ;
      RECT 123.22 427.36 129.66 427.56 ;
      RECT 123.22 428.96 129.66 429.16 ;
      RECT 123.22 430.76 129.66 430.96 ;
      RECT 123.22 432.36 129.66 432.56 ;
      RECT 123.22 434.16 129.66 434.36 ;
      RECT 123.22 435.76 129.66 435.96 ;
      RECT 123.22 437.56 129.66 437.76 ;
      RECT 123.22 439.16 129.66 439.36 ;
      RECT 123.22 440.96 129.66 441.16 ;
      RECT 123.22 442.56 129.66 442.76 ;
      RECT 123.22 444.36 129.66 444.56 ;
      RECT 123.22 445.96 129.66 446.16 ;
      RECT 123.22 447.76 129.66 447.96 ;
      RECT 123.22 449.36 129.66 449.56 ;
      RECT 123.22 451.16 129.66 451.36 ;
      RECT 123.22 452.76 129.66 452.96 ;
      RECT 123.22 454.56 129.66 454.76 ;
      RECT 123.22 456.16 129.66 456.36 ;
      RECT 123.22 457.96 129.66 458.16 ;
      RECT 123.22 459.56 129.66 459.76 ;
      RECT 123.22 461.36 129.66 461.56 ;
      RECT 123.22 462.96 129.66 463.16 ;
      RECT 123.22 464.76 129.66 464.96 ;
      RECT 123.22 466.36 129.66 466.56 ;
      RECT 123.22 468.16 129.66 468.36 ;
      RECT 123.22 469.76 129.66 469.96 ;
      RECT 123.22 471.56 129.66 471.76 ;
      RECT 123.22 473.16 129.66 473.36 ;
      RECT 123.22 474.96 129.66 475.16 ;
      RECT 123.22 476.56 129.66 476.76 ;
      RECT 123.22 478.36 129.66 478.56 ;
      RECT 123.22 479.96 129.66 480.16 ;
      RECT 123.22 481.76 129.66 481.96 ;
      RECT 123.22 483.36 129.66 483.56 ;
      RECT 123.22 485.16 129.66 485.36 ;
      RECT 123.22 486.76 129.66 486.96 ;
      RECT 123.22 488.56 129.66 488.76 ;
      RECT 123.22 490.16 129.66 490.36 ;
      RECT 123.22 491.96 129.66 492.16 ;
      RECT 123.22 493.56 129.66 493.76 ;
      RECT 123.22 495.36 129.66 495.56 ;
      RECT 123.22 496.96 129.66 497.16 ;
      RECT 123.22 498.76 129.66 498.96 ;
      RECT 123.22 500.36 129.66 500.56 ;
      RECT 123.22 502.16 129.66 502.36 ;
      RECT 123.22 503.76 129.66 503.96 ;
      RECT 128.21 13.78 129.23 13.98 ;
      RECT 126.85 30.6 128.93 30.8 ;
      RECT 126.85 51.44 128.93 51.64 ;
      RECT 126.93 12.82 128.01 13.02 ;
      RECT 127.81 16.13 128.01 16.73 ;
      RECT 127.81 62.01 128.01 62.79 ;
      RECT 126.59 12.32 127.61 12.52 ;
      RECT 124.01 15.38 127.61 15.58 ;
      RECT 127.3 37.58 127.61 38.38 ;
      RECT 124.81 510.34 127.61 510.94 ;
      RECT 125.21 6.24 127.19 6.84 ;
      RECT 126.9 37.58 127.1 38.38 ;
      RECT 123.49 30.6 125.57 30.8 ;
      RECT 123.49 51.44 125.57 51.64 ;
      RECT 125.32 37.58 125.52 38.38 ;
      RECT 124.81 37.58 125.12 38.38 ;
      RECT 124.41 16.13 124.61 16.73 ;
      RECT 124.41 62.01 124.61 62.79 ;
      RECT 121.41 510.34 124.21 510.94 ;
      RECT 123.06 506.04 124.02 506.36 ;
      RECT 123.21 71.16 124.01 71.36 ;
      RECT 123.21 74.56 124.01 74.76 ;
      RECT 123.21 77.96 124.01 78.16 ;
      RECT 123.21 81.36 124.01 81.56 ;
      RECT 123.21 84.76 124.01 84.96 ;
      RECT 123.21 88.16 124.01 88.36 ;
      RECT 123.21 91.56 124.01 91.76 ;
      RECT 123.21 94.96 124.01 95.16 ;
      RECT 123.21 98.36 124.01 98.56 ;
      RECT 123.21 101.76 124.01 101.96 ;
      RECT 123.21 105.16 124.01 105.36 ;
      RECT 123.21 108.56 124.01 108.76 ;
      RECT 123.21 111.96 124.01 112.16 ;
      RECT 123.21 115.36 124.01 115.56 ;
      RECT 123.21 118.76 124.01 118.96 ;
      RECT 123.21 122.16 124.01 122.36 ;
      RECT 123.21 125.56 124.01 125.76 ;
      RECT 123.21 128.96 124.01 129.16 ;
      RECT 123.21 132.36 124.01 132.56 ;
      RECT 123.21 135.76 124.01 135.96 ;
      RECT 123.21 139.16 124.01 139.36 ;
      RECT 123.21 142.56 124.01 142.76 ;
      RECT 123.21 145.96 124.01 146.16 ;
      RECT 123.21 149.36 124.01 149.56 ;
      RECT 123.21 152.76 124.01 152.96 ;
      RECT 123.21 156.16 124.01 156.36 ;
      RECT 123.21 159.56 124.01 159.76 ;
      RECT 123.21 162.96 124.01 163.16 ;
      RECT 123.21 166.36 124.01 166.56 ;
      RECT 123.21 169.76 124.01 169.96 ;
      RECT 123.21 173.16 124.01 173.36 ;
      RECT 123.21 176.56 124.01 176.76 ;
      RECT 123.21 179.96 124.01 180.16 ;
      RECT 123.21 183.36 124.01 183.56 ;
      RECT 123.21 186.76 124.01 186.96 ;
      RECT 123.21 190.16 124.01 190.36 ;
      RECT 123.21 193.56 124.01 193.76 ;
      RECT 123.21 196.96 124.01 197.16 ;
      RECT 123.21 200.36 124.01 200.56 ;
      RECT 123.21 203.76 124.01 203.96 ;
      RECT 123.21 207.16 124.01 207.36 ;
      RECT 123.21 210.56 124.01 210.76 ;
      RECT 123.21 213.96 124.01 214.16 ;
      RECT 123.21 217.36 124.01 217.56 ;
      RECT 123.21 220.76 124.01 220.96 ;
      RECT 123.21 224.16 124.01 224.36 ;
      RECT 123.21 227.56 124.01 227.76 ;
      RECT 123.21 230.96 124.01 231.16 ;
      RECT 123.21 234.36 124.01 234.56 ;
      RECT 123.21 237.76 124.01 237.96 ;
      RECT 123.21 241.16 124.01 241.36 ;
      RECT 123.21 244.56 124.01 244.76 ;
      RECT 123.21 247.96 124.01 248.16 ;
      RECT 123.21 251.36 124.01 251.56 ;
      RECT 123.21 254.76 124.01 254.96 ;
      RECT 123.21 258.16 124.01 258.36 ;
      RECT 123.21 261.56 124.01 261.76 ;
      RECT 123.21 264.96 124.01 265.16 ;
      RECT 123.21 268.36 124.01 268.56 ;
      RECT 123.21 271.76 124.01 271.96 ;
      RECT 123.21 275.16 124.01 275.36 ;
      RECT 123.21 278.56 124.01 278.76 ;
      RECT 123.21 281.96 124.01 282.16 ;
      RECT 123.21 285.36 124.01 285.56 ;
      RECT 123.21 288.76 124.01 288.96 ;
      RECT 123.21 292.16 124.01 292.36 ;
      RECT 123.21 295.56 124.01 295.76 ;
      RECT 123.21 298.96 124.01 299.16 ;
      RECT 123.21 302.36 124.01 302.56 ;
      RECT 123.21 305.76 124.01 305.96 ;
      RECT 123.21 309.16 124.01 309.36 ;
      RECT 123.21 312.56 124.01 312.76 ;
      RECT 123.21 315.96 124.01 316.16 ;
      RECT 123.21 319.36 124.01 319.56 ;
      RECT 123.21 322.76 124.01 322.96 ;
      RECT 123.21 326.16 124.01 326.36 ;
      RECT 123.21 329.56 124.01 329.76 ;
      RECT 123.21 332.96 124.01 333.16 ;
      RECT 123.21 336.36 124.01 336.56 ;
      RECT 123.21 339.76 124.01 339.96 ;
      RECT 123.21 343.16 124.01 343.36 ;
      RECT 123.21 346.56 124.01 346.76 ;
      RECT 123.21 349.96 124.01 350.16 ;
      RECT 123.21 353.36 124.01 353.56 ;
      RECT 123.21 356.76 124.01 356.96 ;
      RECT 123.21 360.16 124.01 360.36 ;
      RECT 123.21 363.56 124.01 363.76 ;
      RECT 123.21 366.96 124.01 367.16 ;
      RECT 123.21 370.36 124.01 370.56 ;
      RECT 123.21 373.76 124.01 373.96 ;
      RECT 123.21 377.16 124.01 377.36 ;
      RECT 123.21 380.56 124.01 380.76 ;
      RECT 123.21 383.96 124.01 384.16 ;
      RECT 123.21 387.36 124.01 387.56 ;
      RECT 123.21 390.76 124.01 390.96 ;
      RECT 123.21 394.16 124.01 394.36 ;
      RECT 123.21 397.56 124.01 397.76 ;
      RECT 123.21 400.96 124.01 401.16 ;
      RECT 123.21 404.36 124.01 404.56 ;
      RECT 123.21 407.76 124.01 407.96 ;
      RECT 123.21 411.16 124.01 411.36 ;
      RECT 123.21 414.56 124.01 414.76 ;
      RECT 123.21 417.96 124.01 418.16 ;
      RECT 123.21 421.36 124.01 421.56 ;
      RECT 123.21 424.76 124.01 424.96 ;
      RECT 123.21 428.16 124.01 428.36 ;
      RECT 123.21 431.56 124.01 431.76 ;
      RECT 123.21 434.96 124.01 435.16 ;
      RECT 123.21 438.36 124.01 438.56 ;
      RECT 123.21 441.76 124.01 441.96 ;
      RECT 123.21 445.16 124.01 445.36 ;
      RECT 123.21 448.56 124.01 448.76 ;
      RECT 123.21 451.96 124.01 452.16 ;
      RECT 123.21 455.36 124.01 455.56 ;
      RECT 123.21 458.76 124.01 458.96 ;
      RECT 123.21 462.16 124.01 462.36 ;
      RECT 123.21 465.56 124.01 465.76 ;
      RECT 123.21 468.96 124.01 469.16 ;
      RECT 123.21 472.36 124.01 472.56 ;
      RECT 123.21 475.76 124.01 475.96 ;
      RECT 123.21 479.16 124.01 479.36 ;
      RECT 123.21 482.56 124.01 482.76 ;
      RECT 123.21 485.96 124.01 486.16 ;
      RECT 123.21 489.36 124.01 489.56 ;
      RECT 123.21 492.76 124.01 492.96 ;
      RECT 123.21 496.16 124.01 496.36 ;
      RECT 123.21 499.56 124.01 499.76 ;
      RECT 123.21 502.96 124.01 503.16 ;
      RECT 121.83 6.24 123.81 6.84 ;
      RECT 121.41 13.78 122.43 13.98 ;
      RECT 120.05 30.6 122.13 30.8 ;
      RECT 120.05 51.44 122.13 51.64 ;
      RECT 121.23 66.03 121.71 68.22 ;
      RECT 111.21 35.33 121.61 35.53 ;
      RECT 110.5 70.38 121.58 70.58 ;
      RECT 110.5 83.98 121.58 84.18 ;
      RECT 110.5 97.58 121.58 97.78 ;
      RECT 110.5 111.18 121.58 111.38 ;
      RECT 110.5 124.78 121.58 124.98 ;
      RECT 110.5 138.38 121.58 138.58 ;
      RECT 110.5 151.98 121.58 152.18 ;
      RECT 110.5 165.58 121.58 165.78 ;
      RECT 110.5 179.18 121.58 179.38 ;
      RECT 110.5 192.78 121.58 192.98 ;
      RECT 110.5 206.38 121.58 206.58 ;
      RECT 110.5 219.98 121.58 220.18 ;
      RECT 110.5 233.58 121.58 233.78 ;
      RECT 110.5 247.18 121.58 247.38 ;
      RECT 110.5 260.78 121.58 260.98 ;
      RECT 110.5 274.38 121.58 274.58 ;
      RECT 110.5 287.98 121.58 288.18 ;
      RECT 110.5 301.58 121.58 301.78 ;
      RECT 110.5 315.18 121.58 315.38 ;
      RECT 110.5 328.78 121.58 328.98 ;
      RECT 110.5 342.38 121.58 342.58 ;
      RECT 110.5 355.98 121.58 356.18 ;
      RECT 110.5 369.58 121.58 369.78 ;
      RECT 110.5 383.18 121.58 383.38 ;
      RECT 110.5 396.78 121.58 396.98 ;
      RECT 110.5 410.38 121.58 410.58 ;
      RECT 110.5 423.98 121.58 424.18 ;
      RECT 110.5 437.58 121.58 437.78 ;
      RECT 110.5 451.18 121.58 451.38 ;
      RECT 110.5 464.78 121.58 464.98 ;
      RECT 110.5 478.38 121.58 478.58 ;
      RECT 110.5 491.98 121.58 492.18 ;
      RECT 110.5 75.34 121.48 75.54 ;
      RECT 110.5 77.18 121.48 77.38 ;
      RECT 110.4 82.14 121.48 82.34 ;
      RECT 110.5 88.94 121.48 89.14 ;
      RECT 110.5 90.78 121.48 90.98 ;
      RECT 110.4 95.74 121.48 95.94 ;
      RECT 110.5 102.54 121.48 102.74 ;
      RECT 110.5 104.38 121.48 104.58 ;
      RECT 110.4 109.34 121.48 109.54 ;
      RECT 110.5 116.14 121.48 116.34 ;
      RECT 110.5 117.98 121.48 118.18 ;
      RECT 110.4 122.94 121.48 123.14 ;
      RECT 110.5 129.74 121.48 129.94 ;
      RECT 110.5 131.58 121.48 131.78 ;
      RECT 110.4 136.54 121.48 136.74 ;
      RECT 110.5 143.34 121.48 143.54 ;
      RECT 110.5 145.18 121.48 145.38 ;
      RECT 110.4 150.14 121.48 150.34 ;
      RECT 110.5 156.94 121.48 157.14 ;
      RECT 110.5 158.78 121.48 158.98 ;
      RECT 110.4 163.74 121.48 163.94 ;
      RECT 110.5 170.54 121.48 170.74 ;
      RECT 110.5 172.38 121.48 172.58 ;
      RECT 110.4 177.34 121.48 177.54 ;
      RECT 110.5 184.14 121.48 184.34 ;
      RECT 110.5 185.98 121.48 186.18 ;
      RECT 110.4 190.94 121.48 191.14 ;
      RECT 110.5 197.74 121.48 197.94 ;
      RECT 110.5 199.58 121.48 199.78 ;
      RECT 110.4 204.54 121.48 204.74 ;
      RECT 110.5 211.34 121.48 211.54 ;
      RECT 110.5 213.18 121.48 213.38 ;
      RECT 110.4 218.14 121.48 218.34 ;
      RECT 110.5 224.94 121.48 225.14 ;
      RECT 110.5 226.78 121.48 226.98 ;
      RECT 110.4 231.74 121.48 231.94 ;
      RECT 110.5 238.54 121.48 238.74 ;
      RECT 110.5 240.38 121.48 240.58 ;
      RECT 110.4 245.34 121.48 245.54 ;
      RECT 110.5 252.14 121.48 252.34 ;
      RECT 110.5 253.98 121.48 254.18 ;
      RECT 110.4 258.94 121.48 259.14 ;
      RECT 110.5 265.74 121.48 265.94 ;
      RECT 110.5 267.58 121.48 267.78 ;
      RECT 110.4 272.54 121.48 272.74 ;
      RECT 110.5 279.34 121.48 279.54 ;
      RECT 110.5 281.18 121.48 281.38 ;
      RECT 110.4 286.14 121.48 286.34 ;
      RECT 110.5 292.94 121.48 293.14 ;
      RECT 110.5 294.78 121.48 294.98 ;
      RECT 110.4 299.74 121.48 299.94 ;
      RECT 110.5 306.54 121.48 306.74 ;
      RECT 110.5 308.38 121.48 308.58 ;
      RECT 110.4 313.34 121.48 313.54 ;
      RECT 110.5 320.14 121.48 320.34 ;
      RECT 110.5 321.98 121.48 322.18 ;
      RECT 110.4 326.94 121.48 327.14 ;
      RECT 110.5 333.74 121.48 333.94 ;
      RECT 110.5 335.58 121.48 335.78 ;
      RECT 110.4 340.54 121.48 340.74 ;
      RECT 110.5 347.34 121.48 347.54 ;
      RECT 110.5 349.18 121.48 349.38 ;
      RECT 110.4 354.14 121.48 354.34 ;
      RECT 110.5 360.94 121.48 361.14 ;
      RECT 110.5 362.78 121.48 362.98 ;
      RECT 110.4 367.74 121.48 367.94 ;
      RECT 110.5 374.54 121.48 374.74 ;
      RECT 110.5 376.38 121.48 376.58 ;
      RECT 110.4 381.34 121.48 381.54 ;
      RECT 110.5 388.14 121.48 388.34 ;
      RECT 110.5 389.98 121.48 390.18 ;
      RECT 110.4 394.94 121.48 395.14 ;
      RECT 110.5 401.74 121.48 401.94 ;
      RECT 110.5 403.58 121.48 403.78 ;
      RECT 110.4 408.54 121.48 408.74 ;
      RECT 110.5 415.34 121.48 415.54 ;
      RECT 110.5 417.18 121.48 417.38 ;
      RECT 110.4 422.14 121.48 422.34 ;
      RECT 110.5 428.94 121.48 429.14 ;
      RECT 110.5 430.78 121.48 430.98 ;
      RECT 110.4 435.74 121.48 435.94 ;
      RECT 110.5 442.54 121.48 442.74 ;
      RECT 110.5 444.38 121.48 444.58 ;
      RECT 110.4 449.34 121.48 449.54 ;
      RECT 110.5 456.14 121.48 456.34 ;
      RECT 110.5 457.98 121.48 458.18 ;
      RECT 110.4 462.94 121.48 463.14 ;
      RECT 110.5 469.74 121.48 469.94 ;
      RECT 110.5 471.58 121.48 471.78 ;
      RECT 110.4 476.54 121.48 476.74 ;
      RECT 110.5 483.34 121.48 483.54 ;
      RECT 110.5 485.18 121.48 485.38 ;
      RECT 110.4 490.14 121.48 490.34 ;
      RECT 110.5 496.94 121.48 497.14 ;
      RECT 110.5 498.78 121.48 498.98 ;
      RECT 110.4 503.74 121.48 503.94 ;
      RECT 120.13 12.82 121.21 13.02 ;
      RECT 121.01 16.13 121.21 16.73 ;
      RECT 121.01 62.01 121.21 62.79 ;
      RECT 120.46 66.03 120.94 68.22 ;
      RECT 119.79 12.32 120.81 12.52 ;
      RECT 117.21 34.53 120.81 34.73 ;
      RECT 120.5 37.58 120.81 38.38 ;
      RECT 118.01 506.26 120.81 506.46 ;
      RECT 118.01 507.72 120.81 507.92 ;
      RECT 118.01 510.34 120.81 510.94 ;
      RECT 111.28 71.95 120.8 72.15 ;
      RECT 111.28 85.55 120.8 85.75 ;
      RECT 111.28 99.15 120.8 99.35 ;
      RECT 111.28 112.75 120.8 112.95 ;
      RECT 111.28 126.35 120.8 126.55 ;
      RECT 111.28 139.95 120.8 140.15 ;
      RECT 111.28 153.55 120.8 153.75 ;
      RECT 111.28 167.15 120.8 167.35 ;
      RECT 111.28 180.75 120.8 180.95 ;
      RECT 111.28 194.35 120.8 194.55 ;
      RECT 111.28 207.95 120.8 208.15 ;
      RECT 111.28 221.55 120.8 221.75 ;
      RECT 111.28 235.15 120.8 235.35 ;
      RECT 111.28 248.75 120.8 248.95 ;
      RECT 111.28 262.35 120.8 262.55 ;
      RECT 111.28 275.95 120.8 276.15 ;
      RECT 111.28 289.55 120.8 289.75 ;
      RECT 111.28 303.15 120.8 303.35 ;
      RECT 111.28 316.75 120.8 316.95 ;
      RECT 111.28 330.35 120.8 330.55 ;
      RECT 111.28 343.95 120.8 344.15 ;
      RECT 111.28 357.55 120.8 357.75 ;
      RECT 111.28 371.15 120.8 371.35 ;
      RECT 111.28 384.75 120.8 384.95 ;
      RECT 111.28 398.35 120.8 398.55 ;
      RECT 111.28 411.95 120.8 412.15 ;
      RECT 111.28 425.55 120.8 425.75 ;
      RECT 111.28 439.15 120.8 439.35 ;
      RECT 111.28 452.75 120.8 452.95 ;
      RECT 111.28 466.35 120.8 466.55 ;
      RECT 111.28 479.95 120.8 480.15 ;
      RECT 111.28 493.55 120.8 493.75 ;
      RECT 111.28 73.77 120.7 73.97 ;
      RECT 111.28 78.75 120.7 78.95 ;
      RECT 111.18 80.57 120.7 80.77 ;
      RECT 111.28 87.37 120.7 87.57 ;
      RECT 111.28 92.35 120.7 92.55 ;
      RECT 111.18 94.17 120.7 94.37 ;
      RECT 111.28 100.97 120.7 101.17 ;
      RECT 111.28 105.95 120.7 106.15 ;
      RECT 111.18 107.77 120.7 107.97 ;
      RECT 111.28 114.57 120.7 114.77 ;
      RECT 111.28 119.55 120.7 119.75 ;
      RECT 111.18 121.37 120.7 121.57 ;
      RECT 111.28 128.17 120.7 128.37 ;
      RECT 111.28 133.15 120.7 133.35 ;
      RECT 111.18 134.97 120.7 135.17 ;
      RECT 111.28 141.77 120.7 141.97 ;
      RECT 111.28 146.75 120.7 146.95 ;
      RECT 111.18 148.57 120.7 148.77 ;
      RECT 111.28 155.37 120.7 155.57 ;
      RECT 111.28 160.35 120.7 160.55 ;
      RECT 111.18 162.17 120.7 162.37 ;
      RECT 111.28 168.97 120.7 169.17 ;
      RECT 111.28 173.95 120.7 174.15 ;
      RECT 111.18 175.77 120.7 175.97 ;
      RECT 111.28 182.57 120.7 182.77 ;
      RECT 111.28 187.55 120.7 187.75 ;
      RECT 111.18 189.37 120.7 189.57 ;
      RECT 111.28 196.17 120.7 196.37 ;
      RECT 111.28 201.15 120.7 201.35 ;
      RECT 111.18 202.97 120.7 203.17 ;
      RECT 111.28 209.77 120.7 209.97 ;
      RECT 111.28 214.75 120.7 214.95 ;
      RECT 111.18 216.57 120.7 216.77 ;
      RECT 111.28 223.37 120.7 223.57 ;
      RECT 111.28 228.35 120.7 228.55 ;
      RECT 111.18 230.17 120.7 230.37 ;
      RECT 111.28 236.97 120.7 237.17 ;
      RECT 111.28 241.95 120.7 242.15 ;
      RECT 111.18 243.77 120.7 243.97 ;
      RECT 111.28 250.57 120.7 250.77 ;
      RECT 111.28 255.55 120.7 255.75 ;
      RECT 111.18 257.37 120.7 257.57 ;
      RECT 111.28 264.17 120.7 264.37 ;
      RECT 111.28 269.15 120.7 269.35 ;
      RECT 111.18 270.97 120.7 271.17 ;
      RECT 111.28 277.77 120.7 277.97 ;
      RECT 111.28 282.75 120.7 282.95 ;
      RECT 111.18 284.57 120.7 284.77 ;
      RECT 111.28 291.37 120.7 291.57 ;
      RECT 111.28 296.35 120.7 296.55 ;
      RECT 111.18 298.17 120.7 298.37 ;
      RECT 111.28 304.97 120.7 305.17 ;
      RECT 111.28 309.95 120.7 310.15 ;
      RECT 111.18 311.77 120.7 311.97 ;
      RECT 111.28 318.57 120.7 318.77 ;
      RECT 111.28 323.55 120.7 323.75 ;
      RECT 111.18 325.37 120.7 325.57 ;
      RECT 111.28 332.17 120.7 332.37 ;
      RECT 111.28 337.15 120.7 337.35 ;
      RECT 111.18 338.97 120.7 339.17 ;
      RECT 111.28 345.77 120.7 345.97 ;
      RECT 111.28 350.75 120.7 350.95 ;
      RECT 111.18 352.57 120.7 352.77 ;
      RECT 111.28 359.37 120.7 359.57 ;
      RECT 111.28 364.35 120.7 364.55 ;
      RECT 111.18 366.17 120.7 366.37 ;
      RECT 111.28 372.97 120.7 373.17 ;
      RECT 111.28 377.95 120.7 378.15 ;
      RECT 111.18 379.77 120.7 379.97 ;
      RECT 111.28 386.57 120.7 386.77 ;
      RECT 111.28 391.55 120.7 391.75 ;
      RECT 111.18 393.37 120.7 393.57 ;
      RECT 111.28 400.17 120.7 400.37 ;
      RECT 111.28 405.15 120.7 405.35 ;
      RECT 111.18 406.97 120.7 407.17 ;
      RECT 111.28 413.77 120.7 413.97 ;
      RECT 111.28 418.75 120.7 418.95 ;
      RECT 111.18 420.57 120.7 420.77 ;
      RECT 111.28 427.37 120.7 427.57 ;
      RECT 111.28 432.35 120.7 432.55 ;
      RECT 111.18 434.17 120.7 434.37 ;
      RECT 111.28 440.97 120.7 441.17 ;
      RECT 111.28 445.95 120.7 446.15 ;
      RECT 111.18 447.77 120.7 447.97 ;
      RECT 111.28 454.57 120.7 454.77 ;
      RECT 111.28 459.55 120.7 459.75 ;
      RECT 111.18 461.37 120.7 461.57 ;
      RECT 111.28 468.17 120.7 468.37 ;
      RECT 111.28 473.15 120.7 473.35 ;
      RECT 111.18 474.97 120.7 475.17 ;
      RECT 111.28 481.77 120.7 481.97 ;
      RECT 111.28 486.75 120.7 486.95 ;
      RECT 111.18 488.57 120.7 488.77 ;
      RECT 111.28 495.37 120.7 495.57 ;
      RECT 111.28 500.35 120.7 500.55 ;
      RECT 111.18 502.17 120.7 502.37 ;
      RECT 118.43 6.24 120.39 6.84 ;
      RECT 113.3 32.48 120.3 32.68 ;
      RECT 120.1 37.58 120.3 38.38 ;
      RECT 118.91 69.46 119.91 69.66 ;
      RECT 118.91 72.86 119.91 73.06 ;
      RECT 118.91 76.26 119.91 76.46 ;
      RECT 118.91 79.66 119.91 79.86 ;
      RECT 118.91 83.06 119.91 83.26 ;
      RECT 118.91 86.46 119.91 86.66 ;
      RECT 118.91 89.86 119.91 90.06 ;
      RECT 118.91 93.26 119.91 93.46 ;
      RECT 118.91 96.66 119.91 96.86 ;
      RECT 118.91 100.06 119.91 100.26 ;
      RECT 118.91 103.46 119.91 103.66 ;
      RECT 118.91 106.86 119.91 107.06 ;
      RECT 118.91 110.26 119.91 110.46 ;
      RECT 118.91 113.66 119.91 113.86 ;
      RECT 118.91 117.06 119.91 117.26 ;
      RECT 118.91 120.46 119.91 120.66 ;
      RECT 118.91 123.86 119.91 124.06 ;
      RECT 118.91 127.26 119.91 127.46 ;
      RECT 118.91 130.66 119.91 130.86 ;
      RECT 118.91 134.06 119.91 134.26 ;
      RECT 118.91 137.46 119.91 137.66 ;
      RECT 118.91 140.86 119.91 141.06 ;
      RECT 118.91 144.26 119.91 144.46 ;
      RECT 118.91 147.66 119.91 147.86 ;
      RECT 118.91 151.06 119.91 151.26 ;
      RECT 118.91 154.46 119.91 154.66 ;
      RECT 118.91 157.86 119.91 158.06 ;
      RECT 118.91 161.26 119.91 161.46 ;
      RECT 118.91 164.66 119.91 164.86 ;
      RECT 118.91 168.06 119.91 168.26 ;
      RECT 118.91 171.46 119.91 171.66 ;
      RECT 118.91 174.86 119.91 175.06 ;
      RECT 118.91 178.26 119.91 178.46 ;
      RECT 118.91 181.66 119.91 181.86 ;
      RECT 118.91 185.06 119.91 185.26 ;
      RECT 118.91 188.46 119.91 188.66 ;
      RECT 118.91 191.86 119.91 192.06 ;
      RECT 118.91 195.26 119.91 195.46 ;
      RECT 118.91 198.66 119.91 198.86 ;
      RECT 118.91 202.06 119.91 202.26 ;
      RECT 118.91 205.46 119.91 205.66 ;
      RECT 118.91 208.86 119.91 209.06 ;
      RECT 118.91 212.26 119.91 212.46 ;
      RECT 118.91 215.66 119.91 215.86 ;
      RECT 118.91 219.06 119.91 219.26 ;
      RECT 118.91 222.46 119.91 222.66 ;
      RECT 118.91 225.86 119.91 226.06 ;
      RECT 118.91 229.26 119.91 229.46 ;
      RECT 118.91 232.66 119.91 232.86 ;
      RECT 118.91 236.06 119.91 236.26 ;
      RECT 118.91 239.46 119.91 239.66 ;
      RECT 118.91 242.86 119.91 243.06 ;
      RECT 118.91 246.26 119.91 246.46 ;
      RECT 118.91 249.66 119.91 249.86 ;
      RECT 118.91 253.06 119.91 253.26 ;
      RECT 118.91 256.46 119.91 256.66 ;
      RECT 118.91 259.86 119.91 260.06 ;
      RECT 118.91 263.26 119.91 263.46 ;
      RECT 118.91 266.66 119.91 266.86 ;
      RECT 118.91 270.06 119.91 270.26 ;
      RECT 118.91 273.46 119.91 273.66 ;
      RECT 118.91 276.86 119.91 277.06 ;
      RECT 118.91 280.26 119.91 280.46 ;
      RECT 118.91 283.66 119.91 283.86 ;
      RECT 118.91 287.06 119.91 287.26 ;
      RECT 118.91 290.46 119.91 290.66 ;
      RECT 118.91 293.86 119.91 294.06 ;
      RECT 118.91 297.26 119.91 297.46 ;
      RECT 118.91 300.66 119.91 300.86 ;
      RECT 118.91 304.06 119.91 304.26 ;
      RECT 118.91 307.46 119.91 307.66 ;
      RECT 118.91 310.86 119.91 311.06 ;
      RECT 118.91 314.26 119.91 314.46 ;
      RECT 118.91 317.66 119.91 317.86 ;
      RECT 118.91 321.06 119.91 321.26 ;
      RECT 118.91 324.46 119.91 324.66 ;
      RECT 118.91 327.86 119.91 328.06 ;
      RECT 118.91 331.26 119.91 331.46 ;
      RECT 118.91 334.66 119.91 334.86 ;
      RECT 118.91 338.06 119.91 338.26 ;
      RECT 118.91 341.46 119.91 341.66 ;
      RECT 118.91 344.86 119.91 345.06 ;
      RECT 118.91 348.26 119.91 348.46 ;
      RECT 118.91 351.66 119.91 351.86 ;
      RECT 118.91 355.06 119.91 355.26 ;
      RECT 118.91 358.46 119.91 358.66 ;
      RECT 118.91 361.86 119.91 362.06 ;
      RECT 118.91 365.26 119.91 365.46 ;
      RECT 118.91 368.66 119.91 368.86 ;
      RECT 118.91 372.06 119.91 372.26 ;
      RECT 118.91 375.46 119.91 375.66 ;
      RECT 118.91 378.86 119.91 379.06 ;
      RECT 118.91 382.26 119.91 382.46 ;
      RECT 118.91 385.66 119.91 385.86 ;
      RECT 118.91 389.06 119.91 389.26 ;
      RECT 118.91 392.46 119.91 392.66 ;
      RECT 118.91 395.86 119.91 396.06 ;
      RECT 118.91 399.26 119.91 399.46 ;
      RECT 118.91 402.66 119.91 402.86 ;
      RECT 118.91 406.06 119.91 406.26 ;
      RECT 118.91 409.46 119.91 409.66 ;
      RECT 118.91 412.86 119.91 413.06 ;
      RECT 118.91 416.26 119.91 416.46 ;
      RECT 118.91 419.66 119.91 419.86 ;
      RECT 118.91 423.06 119.91 423.26 ;
      RECT 118.91 426.46 119.91 426.66 ;
      RECT 118.91 429.86 119.91 430.06 ;
      RECT 118.91 433.26 119.91 433.46 ;
      RECT 118.91 436.66 119.91 436.86 ;
      RECT 118.91 440.06 119.91 440.26 ;
      RECT 118.91 443.46 119.91 443.66 ;
      RECT 118.91 446.86 119.91 447.06 ;
      RECT 118.91 450.26 119.91 450.46 ;
      RECT 118.91 453.66 119.91 453.86 ;
      RECT 118.91 457.06 119.91 457.26 ;
      RECT 118.91 460.46 119.91 460.66 ;
      RECT 118.91 463.86 119.91 464.06 ;
      RECT 118.91 467.26 119.91 467.46 ;
      RECT 118.91 470.66 119.91 470.86 ;
      RECT 118.91 474.06 119.91 474.26 ;
      RECT 118.91 477.46 119.91 477.66 ;
      RECT 118.91 480.86 119.91 481.06 ;
      RECT 118.91 484.26 119.91 484.46 ;
      RECT 118.91 487.66 119.91 487.86 ;
      RECT 118.91 491.06 119.91 491.26 ;
      RECT 118.91 494.46 119.91 494.66 ;
      RECT 118.91 497.86 119.91 498.06 ;
      RECT 118.91 501.26 119.91 501.46 ;
      RECT 118.91 504.66 119.91 504.86 ;
      RECT 118.01 12.32 119.03 12.52 ;
      RECT 116.69 30.6 118.77 30.8 ;
      RECT 116.69 51.44 118.77 51.64 ;
      RECT 111.72 34.93 118.72 35.13 ;
      RECT 118.52 37.58 118.72 38.38 ;
      RECT 117.61 12.82 118.69 13.02 ;
      RECT 118.01 37.58 118.32 38.38 ;
      RECT 117.83 66.03 118.31 68.22 ;
      RECT 117.61 16.13 117.81 16.73 ;
      RECT 117.61 62.01 117.81 62.79 ;
      RECT 117.06 66.03 117.54 68.22 ;
      RECT 116.39 13.78 117.41 13.98 ;
      RECT 114.61 510.34 117.41 510.94 ;
      RECT 115.03 6.24 116.99 6.84 ;
      RECT 114.61 34.53 116.8 34.73 ;
      RECT 115.51 69.46 116.51 69.66 ;
      RECT 115.51 76.26 116.51 76.46 ;
      RECT 115.51 83.06 116.51 83.26 ;
      RECT 115.51 89.86 116.51 90.06 ;
      RECT 115.51 96.66 116.51 96.86 ;
      RECT 115.51 103.46 116.51 103.66 ;
      RECT 115.51 110.26 116.51 110.46 ;
      RECT 115.51 117.06 116.51 117.26 ;
      RECT 115.51 123.86 116.51 124.06 ;
      RECT 115.51 130.66 116.51 130.86 ;
      RECT 115.51 137.46 116.51 137.66 ;
      RECT 115.51 144.26 116.51 144.46 ;
      RECT 115.51 151.06 116.51 151.26 ;
      RECT 115.51 157.86 116.51 158.06 ;
      RECT 115.51 164.66 116.51 164.86 ;
      RECT 115.51 171.46 116.51 171.66 ;
      RECT 115.51 178.26 116.51 178.46 ;
      RECT 115.51 185.06 116.51 185.26 ;
      RECT 115.51 191.86 116.51 192.06 ;
      RECT 115.51 198.66 116.51 198.86 ;
      RECT 115.51 205.46 116.51 205.66 ;
      RECT 115.51 212.26 116.51 212.46 ;
      RECT 115.51 219.06 116.51 219.26 ;
      RECT 115.51 225.86 116.51 226.06 ;
      RECT 115.51 232.66 116.51 232.86 ;
      RECT 115.51 239.46 116.51 239.66 ;
      RECT 115.51 246.26 116.51 246.46 ;
      RECT 115.51 253.06 116.51 253.26 ;
      RECT 115.51 259.86 116.51 260.06 ;
      RECT 115.51 266.66 116.51 266.86 ;
      RECT 115.51 273.46 116.51 273.66 ;
      RECT 115.51 280.26 116.51 280.46 ;
      RECT 115.51 287.06 116.51 287.26 ;
      RECT 115.51 293.86 116.51 294.06 ;
      RECT 115.51 300.66 116.51 300.86 ;
      RECT 115.51 307.46 116.51 307.66 ;
      RECT 115.51 314.26 116.51 314.46 ;
      RECT 115.51 321.06 116.51 321.26 ;
      RECT 115.51 327.86 116.51 328.06 ;
      RECT 115.51 334.66 116.51 334.86 ;
      RECT 115.51 341.46 116.51 341.66 ;
      RECT 115.51 348.26 116.51 348.46 ;
      RECT 115.51 355.06 116.51 355.26 ;
      RECT 115.51 361.86 116.51 362.06 ;
      RECT 115.51 368.66 116.51 368.86 ;
      RECT 115.51 375.46 116.51 375.66 ;
      RECT 115.51 382.26 116.51 382.46 ;
      RECT 115.51 389.06 116.51 389.26 ;
      RECT 115.51 395.86 116.51 396.06 ;
      RECT 115.51 402.66 116.51 402.86 ;
      RECT 115.51 409.46 116.51 409.66 ;
      RECT 115.51 416.26 116.51 416.46 ;
      RECT 115.51 423.06 116.51 423.26 ;
      RECT 115.51 429.86 116.51 430.06 ;
      RECT 115.51 436.66 116.51 436.86 ;
      RECT 115.51 443.46 116.51 443.66 ;
      RECT 115.51 450.26 116.51 450.46 ;
      RECT 115.51 457.06 116.51 457.26 ;
      RECT 115.51 463.86 116.51 464.06 ;
      RECT 115.51 470.66 116.51 470.86 ;
      RECT 115.51 477.46 116.51 477.66 ;
      RECT 115.51 484.26 116.51 484.46 ;
      RECT 115.51 491.06 116.51 491.26 ;
      RECT 115.51 497.86 116.51 498.06 ;
      RECT 115.51 504.66 116.51 504.86 ;
      RECT 109.46 70.84 115.79 71.16 ;
      RECT 109.46 74.76 115.79 75.08 ;
      RECT 109.46 77.64 115.79 77.96 ;
      RECT 109.46 81.56 115.79 81.88 ;
      RECT 109.46 84.44 115.79 84.76 ;
      RECT 109.46 88.36 115.79 88.68 ;
      RECT 109.46 91.24 115.79 91.56 ;
      RECT 109.46 95.16 115.79 95.48 ;
      RECT 109.46 98.04 115.79 98.36 ;
      RECT 109.46 101.96 115.79 102.28 ;
      RECT 109.46 104.84 115.79 105.16 ;
      RECT 109.46 108.76 115.79 109.08 ;
      RECT 109.46 111.64 115.79 111.96 ;
      RECT 109.46 115.56 115.79 115.88 ;
      RECT 109.46 118.44 115.79 118.76 ;
      RECT 109.46 122.36 115.79 122.68 ;
      RECT 109.46 125.24 115.79 125.56 ;
      RECT 109.46 129.16 115.79 129.48 ;
      RECT 109.46 132.04 115.79 132.36 ;
      RECT 109.46 135.96 115.79 136.28 ;
      RECT 109.46 138.84 115.79 139.16 ;
      RECT 109.46 142.76 115.79 143.08 ;
      RECT 109.46 145.64 115.79 145.96 ;
      RECT 109.46 149.56 115.79 149.88 ;
      RECT 109.46 152.44 115.79 152.76 ;
      RECT 109.46 156.36 115.79 156.68 ;
      RECT 109.46 159.24 115.79 159.56 ;
      RECT 109.46 163.16 115.79 163.48 ;
      RECT 109.46 166.04 115.79 166.36 ;
      RECT 109.46 169.96 115.79 170.28 ;
      RECT 109.46 172.84 115.79 173.16 ;
      RECT 109.46 176.76 115.79 177.08 ;
      RECT 109.46 179.64 115.79 179.96 ;
      RECT 109.46 183.56 115.79 183.88 ;
      RECT 109.46 186.44 115.79 186.76 ;
      RECT 109.46 190.36 115.79 190.68 ;
      RECT 109.46 193.24 115.79 193.56 ;
      RECT 109.46 197.16 115.79 197.48 ;
      RECT 109.46 200.04 115.79 200.36 ;
      RECT 109.46 203.96 115.79 204.28 ;
      RECT 109.46 206.84 115.79 207.16 ;
      RECT 109.46 210.76 115.79 211.08 ;
      RECT 109.46 213.64 115.79 213.96 ;
      RECT 109.46 217.56 115.79 217.88 ;
      RECT 109.46 220.44 115.79 220.76 ;
      RECT 109.46 224.36 115.79 224.68 ;
      RECT 109.46 227.24 115.79 227.56 ;
      RECT 109.46 231.16 115.79 231.48 ;
      RECT 109.46 234.04 115.79 234.36 ;
      RECT 109.46 237.96 115.79 238.28 ;
      RECT 109.46 240.84 115.79 241.16 ;
      RECT 109.46 244.76 115.79 245.08 ;
      RECT 109.46 247.64 115.79 247.96 ;
      RECT 109.46 251.56 115.79 251.88 ;
      RECT 109.46 254.44 115.79 254.76 ;
      RECT 109.46 258.36 115.79 258.68 ;
      RECT 109.46 261.24 115.79 261.56 ;
      RECT 109.46 265.16 115.79 265.48 ;
      RECT 109.46 268.04 115.79 268.36 ;
      RECT 109.46 271.96 115.79 272.28 ;
      RECT 109.46 274.84 115.79 275.16 ;
      RECT 109.46 278.76 115.79 279.08 ;
      RECT 109.46 281.64 115.79 281.96 ;
      RECT 109.46 285.56 115.79 285.88 ;
      RECT 109.46 288.44 115.79 288.76 ;
      RECT 109.46 292.36 115.79 292.68 ;
      RECT 109.46 295.24 115.79 295.56 ;
      RECT 109.46 299.16 115.79 299.48 ;
      RECT 109.46 302.04 115.79 302.36 ;
      RECT 109.46 305.96 115.79 306.28 ;
      RECT 109.46 308.84 115.79 309.16 ;
      RECT 109.46 312.76 115.79 313.08 ;
      RECT 109.46 315.64 115.79 315.96 ;
      RECT 109.46 319.56 115.79 319.88 ;
      RECT 109.46 322.44 115.79 322.76 ;
      RECT 109.46 326.36 115.79 326.68 ;
      RECT 109.46 329.24 115.79 329.56 ;
      RECT 109.46 333.16 115.79 333.48 ;
      RECT 109.46 336.04 115.79 336.36 ;
      RECT 109.46 339.96 115.79 340.28 ;
      RECT 109.46 342.84 115.79 343.16 ;
      RECT 109.46 346.76 115.79 347.08 ;
      RECT 109.46 349.64 115.79 349.96 ;
      RECT 109.46 353.56 115.79 353.88 ;
      RECT 109.46 356.44 115.79 356.76 ;
      RECT 109.46 360.36 115.79 360.68 ;
      RECT 109.46 363.24 115.79 363.56 ;
      RECT 109.46 367.16 115.79 367.48 ;
      RECT 109.46 370.04 115.79 370.36 ;
      RECT 109.46 373.96 115.79 374.28 ;
      RECT 109.46 376.84 115.79 377.16 ;
      RECT 109.46 380.76 115.79 381.08 ;
      RECT 109.46 383.64 115.79 383.96 ;
      RECT 109.46 387.56 115.79 387.88 ;
      RECT 109.46 390.44 115.79 390.76 ;
      RECT 109.46 394.36 115.79 394.68 ;
      RECT 109.46 397.24 115.79 397.56 ;
      RECT 109.46 401.16 115.79 401.48 ;
      RECT 109.46 404.04 115.79 404.36 ;
      RECT 109.46 407.96 115.79 408.28 ;
      RECT 109.46 410.84 115.79 411.16 ;
      RECT 109.46 414.76 115.79 415.08 ;
      RECT 109.46 417.64 115.79 417.96 ;
      RECT 109.46 421.56 115.79 421.88 ;
      RECT 109.46 424.44 115.79 424.76 ;
      RECT 109.46 428.36 115.79 428.68 ;
      RECT 109.46 431.24 115.79 431.56 ;
      RECT 109.46 435.16 115.79 435.48 ;
      RECT 109.46 438.04 115.79 438.36 ;
      RECT 109.46 441.96 115.79 442.28 ;
      RECT 109.46 444.84 115.79 445.16 ;
      RECT 109.46 448.76 115.79 449.08 ;
      RECT 109.46 451.64 115.79 451.96 ;
      RECT 109.46 455.56 115.79 455.88 ;
      RECT 109.46 458.44 115.79 458.76 ;
      RECT 109.46 462.36 115.79 462.68 ;
      RECT 109.46 465.24 115.79 465.56 ;
      RECT 109.46 469.16 115.79 469.48 ;
      RECT 109.46 472.04 115.79 472.36 ;
      RECT 109.46 475.96 115.79 476.28 ;
      RECT 109.46 478.84 115.79 479.16 ;
      RECT 109.46 482.76 115.79 483.08 ;
      RECT 109.46 485.64 115.79 485.96 ;
      RECT 109.46 489.56 115.79 489.88 ;
      RECT 109.46 492.44 115.79 492.76 ;
      RECT 109.46 496.36 115.79 496.68 ;
      RECT 109.46 499.24 115.79 499.56 ;
      RECT 109.46 503.16 115.79 503.48 ;
      RECT 114.61 13.78 115.63 13.98 ;
      RECT 113.25 30.6 115.33 30.8 ;
      RECT 113.25 51.44 115.33 51.64 ;
      RECT 114.43 66.03 114.91 68.22 ;
      RECT 113.33 12.82 114.41 13.02 ;
      RECT 114.21 16.13 114.41 16.73 ;
      RECT 114.21 62.01 114.41 62.79 ;
      RECT 113.66 66.03 114.14 68.22 ;
      RECT 112.99 12.32 114.01 12.52 ;
      RECT 110.41 15.38 114.01 15.58 ;
      RECT 113.7 37.58 114.01 38.38 ;
      RECT 111.21 510.34 114.01 510.94 ;
      RECT 111.61 6.24 113.59 6.84 ;
      RECT 113.3 37.58 113.5 38.38 ;
      RECT 109.89 30.6 111.97 30.8 ;
      RECT 109.89 51.44 111.97 51.64 ;
      RECT 111.72 37.58 111.92 38.38 ;
      RECT 111.21 37.58 111.52 38.38 ;
      RECT 111.03 66.03 111.51 68.22 ;
      RECT 110.81 16.13 111.01 16.73 ;
      RECT 110.81 62.01 111.01 62.79 ;
      RECT 110.26 66.03 110.74 68.22 ;
      RECT 109.51 510.34 110.61 510.94 ;
      RECT 108.23 6.24 110.21 6.84 ;
      RECT 107.81 510.34 108.91 510.94 ;
      RECT 107.81 13.78 108.83 13.98 ;
      RECT 108.41 68.43 108.81 70.66 ;
      RECT 108.41 70.96 108.81 84.26 ;
      RECT 108.41 84.56 108.81 97.86 ;
      RECT 108.41 98.16 108.81 111.46 ;
      RECT 108.41 111.76 108.81 125.06 ;
      RECT 108.41 125.36 108.81 138.66 ;
      RECT 108.41 138.96 108.81 152.26 ;
      RECT 108.41 152.56 108.81 165.86 ;
      RECT 108.41 166.16 108.81 179.46 ;
      RECT 108.41 179.76 108.81 193.06 ;
      RECT 108.41 193.36 108.81 206.66 ;
      RECT 108.41 206.96 108.81 220.26 ;
      RECT 108.41 220.56 108.81 233.86 ;
      RECT 108.41 234.16 108.81 247.46 ;
      RECT 108.41 247.76 108.81 261.06 ;
      RECT 108.41 261.36 108.81 274.66 ;
      RECT 108.41 274.96 108.81 288.26 ;
      RECT 108.41 288.56 108.81 301.86 ;
      RECT 108.41 302.16 108.81 315.46 ;
      RECT 108.41 315.76 108.81 329.06 ;
      RECT 108.41 329.36 108.81 342.66 ;
      RECT 108.41 342.96 108.81 356.26 ;
      RECT 108.41 356.56 108.81 369.86 ;
      RECT 108.41 370.16 108.81 383.46 ;
      RECT 108.41 383.76 108.81 397.06 ;
      RECT 108.41 397.36 108.81 410.66 ;
      RECT 108.41 410.96 108.81 424.26 ;
      RECT 108.41 424.56 108.81 437.86 ;
      RECT 108.41 438.16 108.81 451.46 ;
      RECT 108.41 451.76 108.81 465.06 ;
      RECT 108.41 465.36 108.81 478.66 ;
      RECT 108.41 478.96 108.81 492.26 ;
      RECT 108.41 492.56 108.81 506.24 ;
      RECT 106.45 30.6 108.53 30.8 ;
      RECT 106.45 51.44 108.53 51.64 ;
      RECT 107.63 66.03 108.11 505.98 ;
      RECT 97.61 35.33 108.01 35.53 ;
      RECT 106.53 12.82 107.61 13.02 ;
      RECT 107.41 16.13 107.61 16.73 ;
      RECT 107.41 62.01 107.61 62.79 ;
      RECT 106.86 66.03 107.34 505.98 ;
      RECT 106.19 12.32 107.21 12.52 ;
      RECT 103.61 34.53 107.21 34.73 ;
      RECT 106.9 37.58 107.21 38.38 ;
      RECT 106.11 510.34 107.21 510.94 ;
      RECT 104.83 6.24 106.79 6.84 ;
      RECT 99.7 32.48 106.7 32.68 ;
      RECT 106.5 37.58 106.7 38.38 ;
      RECT 106.16 68.83 106.56 70.66 ;
      RECT 106.16 71.24 106.56 179.46 ;
      RECT 106.16 180.04 106.56 288.26 ;
      RECT 106.16 288.84 106.56 397.06 ;
      RECT 106.16 397.64 106.56 506.32 ;
      RECT 104.41 12.32 105.43 12.52 ;
      RECT 103.09 30.6 105.17 30.8 ;
      RECT 103.09 51.44 105.17 51.64 ;
      RECT 98.12 34.93 105.12 35.13 ;
      RECT 104.92 37.58 105.12 38.38 ;
      RECT 104.01 12.82 105.09 13.02 ;
      RECT 104.41 37.58 104.72 38.38 ;
      RECT 104.23 66.03 104.71 505.98 ;
      RECT 104.01 16.13 104.21 16.73 ;
      RECT 104.01 62.01 104.21 62.79 ;
      RECT 103.46 66.03 103.94 505.98 ;
      RECT 102.79 13.78 103.81 13.98 ;
      RECT 101.43 6.24 103.39 6.84 ;
      RECT 101.01 34.53 103.2 34.73 ;
      RECT 101.01 13.78 102.03 13.98 ;
      RECT 99.65 30.6 101.73 30.8 ;
      RECT 99.65 51.44 101.73 51.64 ;
      RECT 100.83 66.03 101.31 505.98 ;
      RECT 99.73 12.82 100.81 13.02 ;
      RECT 100.61 16.13 100.81 16.73 ;
      RECT 100.61 62.01 100.81 62.79 ;
      RECT 100.06 66.03 100.54 505.98 ;
      RECT 99.39 12.32 100.41 12.52 ;
      RECT 96.81 15.38 100.41 15.58 ;
      RECT 100.1 37.58 100.41 38.38 ;
      RECT 98.01 6.24 99.99 6.84 ;
      RECT 99.7 37.58 99.9 38.38 ;
      RECT 96.29 30.6 98.37 30.8 ;
      RECT 96.29 51.44 98.37 51.64 ;
      RECT 98.12 37.58 98.32 38.38 ;
      RECT 97.61 37.58 97.92 38.38 ;
      RECT 97.43 66.03 97.91 505.98 ;
      RECT 97.21 16.13 97.41 16.73 ;
      RECT 97.21 62.01 97.41 62.79 ;
      RECT 96.66 66.03 97.14 505.98 ;
      RECT 94.63 6.24 96.61 6.84 ;
      RECT 94.21 13.78 95.23 13.98 ;
      RECT 92.85 30.6 94.93 30.8 ;
      RECT 92.85 51.44 94.93 51.64 ;
      RECT 94.03 66.04 94.51 505.98 ;
      RECT 92.93 12.82 94.01 13.02 ;
      RECT 93.81 16.13 94.01 16.73 ;
      RECT 93.81 62.01 94.01 62.79 ;
      RECT 93.26 66.03 93.74 505.98 ;
      RECT 92.59 12.32 93.61 12.52 ;
      RECT 91.23 6.24 93.19 6.84 ;
      RECT 90.01 32.51 93.11 32.71 ;
      RECT 92.9 37.58 93.1 38.38 ;
      RECT 90.81 12.32 91.83 12.52 ;
      RECT 89.49 30.6 91.57 30.8 ;
      RECT 89.49 51.44 91.57 51.64 ;
      RECT 91.32 37.58 91.52 38.38 ;
      RECT 90.41 12.82 91.49 13.02 ;
      RECT 90.63 66.04 91.11 505.98 ;
      RECT 90.41 16.13 90.61 16.73 ;
      RECT 90.41 62.01 90.61 62.79 ;
      RECT 89.86 66.03 90.34 505.98 ;
      RECT 89.19 13.78 90.21 13.98 ;
      RECT 88.81 6.24 89.79 6.84 ;
      RECT 87.21 6.24 88.01 6.64 ;
      RECT 6.83 19.01 88.01 19.81 ;
      RECT 8.21 52.04 88.01 52.84 ;
      RECT 6.24 57.02 87.41 58.02 ;
      RECT 6.24 31.13 87.11 32.13 ;
      RECT 86.91 69.4 87.11 70.2 ;
      RECT 86.91 70.4 87.11 71.16 ;
      RECT 86.91 71.36 87.11 72.12 ;
      RECT 86.91 72.32 87.11 73.6 ;
      RECT 86.91 73.8 87.11 74.56 ;
      RECT 86.91 74.76 87.11 75.52 ;
      RECT 86.91 75.72 87.11 77 ;
      RECT 86.91 77.2 87.11 77.96 ;
      RECT 86.91 78.16 87.11 78.92 ;
      RECT 86.91 79.12 87.11 80.4 ;
      RECT 86.91 80.6 87.11 81.36 ;
      RECT 86.91 81.56 87.11 82.32 ;
      RECT 86.91 82.52 87.11 83.8 ;
      RECT 86.91 84 87.11 84.76 ;
      RECT 86.91 84.96 87.11 85.72 ;
      RECT 86.91 85.92 87.11 87.2 ;
      RECT 86.91 87.4 87.11 88.16 ;
      RECT 86.91 88.36 87.11 89.12 ;
      RECT 86.91 89.32 87.11 90.6 ;
      RECT 86.91 90.8 87.11 91.56 ;
      RECT 86.91 91.76 87.11 92.52 ;
      RECT 86.91 92.72 87.11 94 ;
      RECT 86.91 94.2 87.11 94.96 ;
      RECT 86.91 95.16 87.11 95.92 ;
      RECT 86.91 96.12 87.11 97.4 ;
      RECT 86.91 97.6 87.11 98.36 ;
      RECT 86.91 98.56 87.11 99.32 ;
      RECT 86.91 99.52 87.11 100.8 ;
      RECT 86.91 101 87.11 101.76 ;
      RECT 86.91 101.96 87.11 102.72 ;
      RECT 86.91 102.92 87.11 104.2 ;
      RECT 86.91 104.4 87.11 105.16 ;
      RECT 86.91 105.36 87.11 106.12 ;
      RECT 86.91 106.32 87.11 107.6 ;
      RECT 86.91 107.8 87.11 108.56 ;
      RECT 86.91 108.76 87.11 109.52 ;
      RECT 86.91 109.72 87.11 111 ;
      RECT 86.91 111.2 87.11 111.96 ;
      RECT 86.91 112.16 87.11 112.92 ;
      RECT 86.91 113.12 87.11 114.4 ;
      RECT 86.91 114.6 87.11 115.36 ;
      RECT 86.91 115.56 87.11 116.32 ;
      RECT 86.91 116.52 87.11 117.8 ;
      RECT 86.91 118 87.11 118.76 ;
      RECT 86.91 118.96 87.11 119.72 ;
      RECT 86.91 119.92 87.11 121.2 ;
      RECT 86.91 121.4 87.11 122.16 ;
      RECT 86.91 122.36 87.11 123.12 ;
      RECT 86.91 123.32 87.11 124.6 ;
      RECT 86.91 124.8 87.11 125.56 ;
      RECT 86.91 125.76 87.11 126.52 ;
      RECT 86.91 126.72 87.11 128 ;
      RECT 86.91 128.2 87.11 128.96 ;
      RECT 86.91 129.16 87.11 129.92 ;
      RECT 86.91 130.12 87.11 131.4 ;
      RECT 86.91 131.6 87.11 132.36 ;
      RECT 86.91 132.56 87.11 133.32 ;
      RECT 86.91 133.52 87.11 134.8 ;
      RECT 86.91 135 87.11 135.76 ;
      RECT 86.91 135.96 87.11 136.72 ;
      RECT 86.91 136.92 87.11 138.2 ;
      RECT 86.91 138.4 87.11 139.16 ;
      RECT 86.91 139.36 87.11 140.12 ;
      RECT 86.91 140.32 87.11 141.6 ;
      RECT 86.91 141.8 87.11 142.56 ;
      RECT 86.91 142.76 87.11 143.52 ;
      RECT 86.91 143.72 87.11 145 ;
      RECT 86.91 145.2 87.11 145.96 ;
      RECT 86.91 146.16 87.11 146.92 ;
      RECT 86.91 147.12 87.11 148.4 ;
      RECT 86.91 148.6 87.11 149.36 ;
      RECT 86.91 149.56 87.11 150.32 ;
      RECT 86.91 150.52 87.11 151.8 ;
      RECT 86.91 152 87.11 152.76 ;
      RECT 86.91 152.96 87.11 153.72 ;
      RECT 86.91 153.92 87.11 155.2 ;
      RECT 86.91 155.4 87.11 156.16 ;
      RECT 86.91 156.36 87.11 157.12 ;
      RECT 86.91 157.32 87.11 158.6 ;
      RECT 86.91 158.8 87.11 159.56 ;
      RECT 86.91 159.76 87.11 160.52 ;
      RECT 86.91 160.72 87.11 162 ;
      RECT 86.91 162.2 87.11 162.96 ;
      RECT 86.91 163.16 87.11 163.92 ;
      RECT 86.91 164.12 87.11 165.4 ;
      RECT 86.91 165.6 87.11 166.36 ;
      RECT 86.91 166.56 87.11 167.32 ;
      RECT 86.91 167.52 87.11 168.8 ;
      RECT 86.91 169 87.11 169.76 ;
      RECT 86.91 169.96 87.11 170.72 ;
      RECT 86.91 170.92 87.11 172.2 ;
      RECT 86.91 172.4 87.11 173.16 ;
      RECT 86.91 173.36 87.11 174.12 ;
      RECT 86.91 174.32 87.11 175.6 ;
      RECT 86.91 175.8 87.11 176.56 ;
      RECT 86.91 176.76 87.11 177.52 ;
      RECT 86.91 177.72 87.11 179 ;
      RECT 86.91 179.2 87.11 179.96 ;
      RECT 86.91 180.16 87.11 180.92 ;
      RECT 86.91 181.12 87.11 182.4 ;
      RECT 86.91 182.6 87.11 183.36 ;
      RECT 86.91 183.56 87.11 184.32 ;
      RECT 86.91 184.52 87.11 185.8 ;
      RECT 86.91 186 87.11 186.76 ;
      RECT 86.91 186.96 87.11 187.72 ;
      RECT 86.91 187.92 87.11 189.2 ;
      RECT 86.91 189.4 87.11 190.16 ;
      RECT 86.91 190.36 87.11 191.12 ;
      RECT 86.91 191.32 87.11 192.6 ;
      RECT 86.91 192.8 87.11 193.56 ;
      RECT 86.91 193.76 87.11 194.52 ;
      RECT 86.91 194.72 87.11 196 ;
      RECT 86.91 196.2 87.11 196.96 ;
      RECT 86.91 197.16 87.11 197.92 ;
      RECT 86.91 198.12 87.11 199.4 ;
      RECT 86.91 199.6 87.11 200.36 ;
      RECT 86.91 200.56 87.11 201.32 ;
      RECT 86.91 201.52 87.11 202.8 ;
      RECT 86.91 203 87.11 203.76 ;
      RECT 86.91 203.96 87.11 204.72 ;
      RECT 86.91 204.92 87.11 206.2 ;
      RECT 86.91 206.4 87.11 207.16 ;
      RECT 86.91 207.36 87.11 208.12 ;
      RECT 86.91 208.32 87.11 209.6 ;
      RECT 86.91 209.8 87.11 210.56 ;
      RECT 86.91 210.76 87.11 211.52 ;
      RECT 86.91 211.72 87.11 213 ;
      RECT 86.91 213.2 87.11 213.96 ;
      RECT 86.91 214.16 87.11 214.92 ;
      RECT 86.91 215.12 87.11 216.4 ;
      RECT 86.91 216.6 87.11 217.36 ;
      RECT 86.91 217.56 87.11 218.32 ;
      RECT 86.91 218.52 87.11 219.8 ;
      RECT 86.91 220 87.11 220.76 ;
      RECT 86.91 220.96 87.11 221.72 ;
      RECT 86.91 221.92 87.11 223.2 ;
      RECT 86.91 223.4 87.11 224.16 ;
      RECT 86.91 224.36 87.11 225.12 ;
      RECT 86.91 225.32 87.11 226.6 ;
      RECT 86.91 226.8 87.11 227.56 ;
      RECT 86.91 227.76 87.11 228.52 ;
      RECT 86.91 228.72 87.11 230 ;
      RECT 86.91 230.2 87.11 230.96 ;
      RECT 86.91 231.16 87.11 231.92 ;
      RECT 86.91 232.12 87.11 233.4 ;
      RECT 86.91 233.6 87.11 234.36 ;
      RECT 86.91 234.56 87.11 235.32 ;
      RECT 86.91 235.52 87.11 236.8 ;
      RECT 86.91 237 87.11 237.76 ;
      RECT 86.91 237.96 87.11 238.72 ;
      RECT 86.91 238.92 87.11 240.2 ;
      RECT 86.91 240.4 87.11 241.16 ;
      RECT 86.91 241.36 87.11 242.12 ;
      RECT 86.91 242.32 87.11 243.6 ;
      RECT 86.91 243.8 87.11 244.56 ;
      RECT 86.91 244.76 87.11 245.52 ;
      RECT 86.91 245.72 87.11 247 ;
      RECT 86.91 247.2 87.11 247.96 ;
      RECT 86.91 248.16 87.11 248.92 ;
      RECT 86.91 249.12 87.11 250.4 ;
      RECT 86.91 250.6 87.11 251.36 ;
      RECT 86.91 251.56 87.11 252.32 ;
      RECT 86.91 252.52 87.11 253.8 ;
      RECT 86.91 254 87.11 254.76 ;
      RECT 86.91 254.96 87.11 255.72 ;
      RECT 86.91 255.92 87.11 257.2 ;
      RECT 86.91 257.4 87.11 258.16 ;
      RECT 86.91 258.36 87.11 259.12 ;
      RECT 86.91 259.32 87.11 260.6 ;
      RECT 86.91 260.8 87.11 261.56 ;
      RECT 86.91 261.76 87.11 262.52 ;
      RECT 86.91 262.72 87.11 264 ;
      RECT 86.91 264.2 87.11 264.96 ;
      RECT 86.91 265.16 87.11 265.92 ;
      RECT 86.91 266.12 87.11 267.4 ;
      RECT 86.91 267.6 87.11 268.36 ;
      RECT 86.91 268.56 87.11 269.32 ;
      RECT 86.91 269.52 87.11 270.8 ;
      RECT 86.91 271 87.11 271.76 ;
      RECT 86.91 271.96 87.11 272.72 ;
      RECT 86.91 272.92 87.11 274.2 ;
      RECT 86.91 274.4 87.11 275.16 ;
      RECT 86.91 275.36 87.11 276.12 ;
      RECT 86.91 276.32 87.11 277.6 ;
      RECT 86.91 277.8 87.11 278.56 ;
      RECT 86.91 278.76 87.11 279.52 ;
      RECT 86.91 279.72 87.11 281 ;
      RECT 86.91 281.2 87.11 281.96 ;
      RECT 86.91 282.16 87.11 282.92 ;
      RECT 86.91 283.12 87.11 284.4 ;
      RECT 86.91 284.6 87.11 285.36 ;
      RECT 86.91 285.56 87.11 286.32 ;
      RECT 86.91 286.52 87.11 287.8 ;
      RECT 86.91 288 87.11 288.76 ;
      RECT 86.91 288.96 87.11 289.72 ;
      RECT 86.91 289.92 87.11 291.2 ;
      RECT 86.91 291.4 87.11 292.16 ;
      RECT 86.91 292.36 87.11 293.12 ;
      RECT 86.91 293.32 87.11 294.6 ;
      RECT 86.91 294.8 87.11 295.56 ;
      RECT 86.91 295.76 87.11 296.52 ;
      RECT 86.91 296.72 87.11 298 ;
      RECT 86.91 298.2 87.11 298.96 ;
      RECT 86.91 299.16 87.11 299.92 ;
      RECT 86.91 300.12 87.11 301.4 ;
      RECT 86.91 301.6 87.11 302.36 ;
      RECT 86.91 302.56 87.11 303.32 ;
      RECT 86.91 303.52 87.11 304.8 ;
      RECT 86.91 305 87.11 305.76 ;
      RECT 86.91 305.96 87.11 306.72 ;
      RECT 86.91 306.92 87.11 308.2 ;
      RECT 86.91 308.4 87.11 309.16 ;
      RECT 86.91 309.36 87.11 310.12 ;
      RECT 86.91 310.32 87.11 311.6 ;
      RECT 86.91 311.8 87.11 312.56 ;
      RECT 86.91 312.76 87.11 313.52 ;
      RECT 86.91 313.72 87.11 315 ;
      RECT 86.91 315.2 87.11 315.96 ;
      RECT 86.91 316.16 87.11 316.92 ;
      RECT 86.91 317.12 87.11 318.4 ;
      RECT 86.91 318.6 87.11 319.36 ;
      RECT 86.91 319.56 87.11 320.32 ;
      RECT 86.91 320.52 87.11 321.8 ;
      RECT 86.91 322 87.11 322.76 ;
      RECT 86.91 322.96 87.11 323.72 ;
      RECT 86.91 323.92 87.11 325.2 ;
      RECT 86.91 325.4 87.11 326.16 ;
      RECT 86.91 326.36 87.11 327.12 ;
      RECT 86.91 327.32 87.11 328.6 ;
      RECT 86.91 328.8 87.11 329.56 ;
      RECT 86.91 329.76 87.11 330.52 ;
      RECT 86.91 330.72 87.11 332 ;
      RECT 86.91 332.2 87.11 332.96 ;
      RECT 86.91 333.16 87.11 333.92 ;
      RECT 86.91 334.12 87.11 335.4 ;
      RECT 86.91 335.6 87.11 336.36 ;
      RECT 86.91 336.56 87.11 337.32 ;
      RECT 86.91 337.52 87.11 338.8 ;
      RECT 86.91 339 87.11 339.76 ;
      RECT 86.91 339.96 87.11 340.72 ;
      RECT 86.91 340.92 87.11 342.2 ;
      RECT 86.91 342.4 87.11 343.16 ;
      RECT 86.91 343.36 87.11 344.12 ;
      RECT 86.91 344.32 87.11 345.6 ;
      RECT 86.91 345.8 87.11 346.56 ;
      RECT 86.91 346.76 87.11 347.52 ;
      RECT 86.91 347.72 87.11 349 ;
      RECT 86.91 349.2 87.11 349.96 ;
      RECT 86.91 350.16 87.11 350.92 ;
      RECT 86.91 351.12 87.11 352.4 ;
      RECT 86.91 352.6 87.11 353.36 ;
      RECT 86.91 353.56 87.11 354.32 ;
      RECT 86.91 354.52 87.11 355.8 ;
      RECT 86.91 356 87.11 356.76 ;
      RECT 86.91 356.96 87.11 357.72 ;
      RECT 86.91 357.92 87.11 359.2 ;
      RECT 86.91 359.4 87.11 360.16 ;
      RECT 86.91 360.36 87.11 361.12 ;
      RECT 86.91 361.32 87.11 362.6 ;
      RECT 86.91 362.8 87.11 363.56 ;
      RECT 86.91 363.76 87.11 364.52 ;
      RECT 86.91 364.72 87.11 366 ;
      RECT 86.91 366.2 87.11 366.96 ;
      RECT 86.91 367.16 87.11 367.92 ;
      RECT 86.91 368.12 87.11 369.4 ;
      RECT 86.91 369.6 87.11 370.36 ;
      RECT 86.91 370.56 87.11 371.32 ;
      RECT 86.91 371.52 87.11 372.8 ;
      RECT 86.91 373 87.11 373.76 ;
      RECT 86.91 373.96 87.11 374.72 ;
      RECT 86.91 374.92 87.11 376.2 ;
      RECT 86.91 376.4 87.11 377.16 ;
      RECT 86.91 377.36 87.11 378.12 ;
      RECT 86.91 378.32 87.11 379.6 ;
      RECT 86.91 379.8 87.11 380.56 ;
      RECT 86.91 380.76 87.11 381.52 ;
      RECT 86.91 381.72 87.11 383 ;
      RECT 86.91 383.2 87.11 383.96 ;
      RECT 86.91 384.16 87.11 384.92 ;
      RECT 86.91 385.12 87.11 386.4 ;
      RECT 86.91 386.6 87.11 387.36 ;
      RECT 86.91 387.56 87.11 388.32 ;
      RECT 86.91 388.52 87.11 389.8 ;
      RECT 86.91 390 87.11 390.76 ;
      RECT 86.91 390.96 87.11 391.72 ;
      RECT 86.91 391.92 87.11 393.2 ;
      RECT 86.91 393.4 87.11 394.16 ;
      RECT 86.91 394.36 87.11 395.12 ;
      RECT 86.91 395.32 87.11 396.6 ;
      RECT 86.91 396.8 87.11 397.56 ;
      RECT 86.91 397.76 87.11 398.52 ;
      RECT 86.91 398.72 87.11 400 ;
      RECT 86.91 400.2 87.11 400.96 ;
      RECT 86.91 401.16 87.11 401.92 ;
      RECT 86.91 402.12 87.11 403.4 ;
      RECT 86.91 403.6 87.11 404.36 ;
      RECT 86.91 404.56 87.11 405.32 ;
      RECT 86.91 405.52 87.11 406.8 ;
      RECT 86.91 407 87.11 407.76 ;
      RECT 86.91 407.96 87.11 408.72 ;
      RECT 86.91 408.92 87.11 410.2 ;
      RECT 86.91 410.4 87.11 411.16 ;
      RECT 86.91 411.36 87.11 412.12 ;
      RECT 86.91 412.32 87.11 413.6 ;
      RECT 86.91 413.8 87.11 414.56 ;
      RECT 86.91 414.76 87.11 415.52 ;
      RECT 86.91 415.72 87.11 417 ;
      RECT 86.91 417.2 87.11 417.96 ;
      RECT 86.91 418.16 87.11 418.92 ;
      RECT 86.91 419.12 87.11 420.4 ;
      RECT 86.91 420.6 87.11 421.36 ;
      RECT 86.91 421.56 87.11 422.32 ;
      RECT 86.91 422.52 87.11 423.8 ;
      RECT 86.91 424 87.11 424.76 ;
      RECT 86.91 424.96 87.11 425.72 ;
      RECT 86.91 425.92 87.11 427.2 ;
      RECT 86.91 427.4 87.11 428.16 ;
      RECT 86.91 428.36 87.11 429.12 ;
      RECT 86.91 429.32 87.11 430.6 ;
      RECT 86.91 430.8 87.11 431.56 ;
      RECT 86.91 431.76 87.11 432.52 ;
      RECT 86.91 432.72 87.11 434 ;
      RECT 86.91 434.2 87.11 434.96 ;
      RECT 86.91 435.16 87.11 435.92 ;
      RECT 86.91 436.12 87.11 437.4 ;
      RECT 86.91 437.6 87.11 438.36 ;
      RECT 86.91 438.56 87.11 439.32 ;
      RECT 86.91 439.52 87.11 440.8 ;
      RECT 86.91 441 87.11 441.76 ;
      RECT 86.91 441.96 87.11 442.72 ;
      RECT 86.91 442.92 87.11 444.2 ;
      RECT 86.91 444.4 87.11 445.16 ;
      RECT 86.91 445.36 87.11 446.12 ;
      RECT 86.91 446.32 87.11 447.6 ;
      RECT 86.91 447.8 87.11 448.56 ;
      RECT 86.91 448.76 87.11 449.52 ;
      RECT 86.91 449.72 87.11 451 ;
      RECT 86.91 451.2 87.11 451.96 ;
      RECT 86.91 452.16 87.11 452.92 ;
      RECT 86.91 453.12 87.11 454.4 ;
      RECT 86.91 454.6 87.11 455.36 ;
      RECT 86.91 455.56 87.11 456.32 ;
      RECT 86.91 456.52 87.11 457.8 ;
      RECT 86.91 458 87.11 458.76 ;
      RECT 86.91 458.96 87.11 459.72 ;
      RECT 86.91 459.92 87.11 461.2 ;
      RECT 86.91 461.4 87.11 462.16 ;
      RECT 86.91 462.36 87.11 463.12 ;
      RECT 86.91 463.32 87.11 464.6 ;
      RECT 86.91 464.8 87.11 465.56 ;
      RECT 86.91 465.76 87.11 466.52 ;
      RECT 86.91 466.72 87.11 468 ;
      RECT 86.91 468.2 87.11 468.96 ;
      RECT 86.91 469.16 87.11 469.92 ;
      RECT 86.91 470.12 87.11 471.4 ;
      RECT 86.91 471.6 87.11 472.36 ;
      RECT 86.91 472.56 87.11 473.32 ;
      RECT 86.91 473.52 87.11 474.8 ;
      RECT 86.91 475 87.11 475.76 ;
      RECT 86.91 475.96 87.11 476.72 ;
      RECT 86.91 476.92 87.11 478.2 ;
      RECT 86.91 478.4 87.11 479.16 ;
      RECT 86.91 479.36 87.11 480.12 ;
      RECT 86.91 480.32 87.11 481.6 ;
      RECT 86.91 481.8 87.11 482.56 ;
      RECT 86.91 482.76 87.11 483.52 ;
      RECT 86.91 483.72 87.11 485 ;
      RECT 86.91 485.2 87.11 485.96 ;
      RECT 86.91 486.16 87.11 486.92 ;
      RECT 86.91 487.12 87.11 488.4 ;
      RECT 86.91 488.6 87.11 489.36 ;
      RECT 86.91 489.56 87.11 490.32 ;
      RECT 86.91 490.52 87.11 491.8 ;
      RECT 86.91 492 87.11 492.76 ;
      RECT 86.91 492.96 87.11 493.72 ;
      RECT 86.91 493.92 87.11 495.2 ;
      RECT 86.91 495.4 87.11 496.16 ;
      RECT 86.91 496.36 87.11 497.12 ;
      RECT 86.91 497.32 87.11 498.6 ;
      RECT 86.91 498.8 87.11 499.56 ;
      RECT 86.91 499.76 87.11 500.52 ;
      RECT 86.91 500.72 87.11 502 ;
      RECT 86.91 502.2 87.11 502.96 ;
      RECT 86.91 503.16 87.11 503.92 ;
      RECT 86.91 504.12 87.11 506.44 ;
      RECT 86.91 506.64 87.11 507.4 ;
      RECT 86.91 507.6 87.11 508.36 ;
      RECT 86.91 508.56 87.11 510 ;
      RECT 85.41 6.24 86.71 6.84 ;
      RECT 86.11 505.38 86.31 510.01 ;
      RECT 85.51 35.31 86.11 35.51 ;
      RECT 85.59 30.13 85.91 30.73 ;
      RECT 85.59 42.75 85.91 43.35 ;
      RECT 77.51 28.15 85.71 28.75 ;
      RECT 84.91 59.37 85.55 59.97 ;
      RECT 66.61 35.75 85.51 35.95 ;
      RECT 66.61 37.21 85.51 37.41 ;
      RECT 85.31 63.99 85.51 505.18 ;
      RECT 85.31 505.38 85.51 510.01 ;
      RECT 66.61 34.65 85.31 34.85 ;
      RECT 84.91 505.38 85.11 510.01 ;
      RECT 83.03 6.24 85.01 6.84 ;
      RECT 84.31 35.31 84.91 35.51 ;
      RECT 84.51 30.13 84.83 30.73 ;
      RECT 84.51 42.75 84.83 43.35 ;
      RECT 84.11 505.38 84.31 510.01 ;
      RECT 83.71 505.38 83.91 510.01 ;
      RECT 83.11 35.31 83.71 35.51 ;
      RECT 83.19 30.13 83.51 30.73 ;
      RECT 83.19 42.75 83.51 43.35 ;
      RECT 83.31 65.96 83.51 510.01 ;
      RECT 82.47 59.37 83.11 59.97 ;
      RECT 82.91 505.38 83.11 510.01 ;
      RECT 82.51 63.99 82.71 505.18 ;
      RECT 82.51 505.38 82.71 510.01 ;
      RECT 80.63 6.24 82.61 6.84 ;
      RECT 81.91 35.31 82.51 35.51 ;
      RECT 82.11 30.13 82.43 30.73 ;
      RECT 82.11 42.75 82.43 43.35 ;
      RECT 80.91 15.51 82.31 15.71 ;
      RECT 82.11 65.96 82.31 510.01 ;
      RECT 81.71 505.38 81.91 510.01 ;
      RECT 81.31 505.38 81.51 510.01 ;
      RECT 80.71 35.31 81.31 35.51 ;
      RECT 80.79 30.13 81.11 30.73 ;
      RECT 80.79 42.75 81.11 43.35 ;
      RECT 80.11 59.37 80.75 59.97 ;
      RECT 80.51 63.99 80.71 505.18 ;
      RECT 80.51 505.38 80.71 510.01 ;
      RECT 80.11 505.38 80.31 510.01 ;
      RECT 78.23 6.24 80.21 6.84 ;
      RECT 79.51 35.31 80.11 35.51 ;
      RECT 79.71 30.13 80.03 30.73 ;
      RECT 79.71 42.75 80.03 43.35 ;
      RECT 79.31 505.38 79.51 510.01 ;
      RECT 78.91 505.38 79.11 510.01 ;
      RECT 78.31 35.31 78.91 35.51 ;
      RECT 78.39 30.13 78.71 30.73 ;
      RECT 78.39 42.75 78.71 43.35 ;
      RECT 78.51 65.96 78.71 510.01 ;
      RECT 77.67 59.37 78.31 59.97 ;
      RECT 78.11 505.38 78.31 510.01 ;
      RECT 77.71 63.99 77.91 505.18 ;
      RECT 77.71 505.38 77.91 510.01 ;
      RECT 75.81 6.24 77.81 6.84 ;
      RECT 77.11 35.31 77.71 35.51 ;
      RECT 77.31 30.13 77.63 30.73 ;
      RECT 77.31 42.75 77.63 43.35 ;
      RECT 77.31 65.96 77.51 510.01 ;
      RECT 76.65 12.98 77.25 13.18 ;
      RECT 76.91 505.38 77.11 510.01 ;
      RECT 76.51 505.38 76.71 510.01 ;
      RECT 75.55 8.94 76.51 9.14 ;
      RECT 75.91 35.31 76.51 35.51 ;
      RECT 72.05 13.78 76.41 13.98 ;
      RECT 75.99 30.13 76.31 30.73 ;
      RECT 75.99 42.75 76.31 43.35 ;
      RECT 75.96 28.03 76.16 28.77 ;
      RECT 68.01 21.31 76.01 21.51 ;
      RECT 74.05 20.61 76 21.01 ;
      RECT 75.31 59.37 75.95 59.97 ;
      RECT 75.71 63.99 75.91 505.18 ;
      RECT 75.71 505.38 75.91 510.01 ;
      RECT 74.72 16.58 75.76 16.78 ;
      RECT 68.26 27.51 75.76 27.71 ;
      RECT 68.26 27.91 75.76 28.11 ;
      RECT 75.31 505.38 75.51 510.01 ;
      RECT 73.44 6.24 75.41 6.84 ;
      RECT 74.71 35.31 75.31 35.51 ;
      RECT 68.73 22.31 75.29 22.51 ;
      RECT 74.91 30.13 75.23 30.73 ;
      RECT 74.91 42.75 75.23 43.35 ;
      RECT 68.97 9.98 75.09 10.18 ;
      RECT 73.97 23.11 75.01 23.31 ;
      RECT 67.71 13.38 74.89 13.58 ;
      RECT 74.11 28.72 74.71 28.92 ;
      RECT 74.51 505.38 74.71 510.01 ;
      RECT 73.97 8.94 74.57 9.14 ;
      RECT 74.11 505.38 74.31 510.01 ;
      RECT 73.2 15.39 74.28 15.59 ;
      RECT 69.85 28.31 74.17 28.51 ;
      RECT 73.51 35.31 74.11 35.51 ;
      RECT 73.41 12.98 74.01 13.18 ;
      RECT 73.59 30.13 73.91 30.73 ;
      RECT 73.59 42.75 73.91 43.35 ;
      RECT 73.71 65.96 73.91 510.01 ;
      RECT 73.55 24.3 73.75 25.07 ;
      RECT 70.35 20.79 73.67 20.99 ;
      RECT 72.87 59.37 73.51 59.97 ;
      RECT 73.31 505.38 73.51 510.01 ;
      RECT 71.41 8.94 73.13 9.14 ;
      RECT 72.91 63.99 73.11 505.18 ;
      RECT 72.91 505.38 73.11 510.01 ;
      RECT 71.51 6.24 73.01 6.84 ;
      RECT 72.31 35.31 72.91 35.51 ;
      RECT 72.51 30.13 72.83 30.73 ;
      RECT 72.51 42.75 72.83 43.35 ;
      RECT 72.51 65.96 72.71 510.01 ;
      RECT 71.61 15.38 72.61 15.72 ;
      RECT 71.45 20.38 72.57 20.58 ;
      RECT 72.11 505.38 72.31 510.01 ;
      RECT 71.71 505.38 71.91 510.01 ;
      RECT 71.11 35.31 71.71 35.51 ;
      RECT 71.19 30.13 71.51 30.73 ;
      RECT 71.19 42.75 71.51 43.35 ;
      RECT 67.61 16.5 71.47 16.7 ;
      RECT 69.61 15.38 71.29 15.58 ;
      RECT 70.61 8.94 71.21 9.14 ;
      RECT 70.51 59.37 71.15 59.97 ;
      RECT 70.91 63.99 71.11 505.18 ;
      RECT 70.91 505.38 71.11 510.01 ;
      RECT 70.51 505.38 70.71 510.01 ;
      RECT 69.09 12.58 70.51 12.78 ;
      RECT 69.91 35.31 70.51 35.51 ;
      RECT 70.27 24.3 70.47 25.07 ;
      RECT 70.11 30.13 70.43 30.73 ;
      RECT 70.11 42.75 70.43 43.35 ;
      RECT 69.61 18.61 70.21 18.81 ;
      RECT 69.11 6.24 70.11 6.84 ;
      RECT 69.01 23.11 70.05 23.31 ;
      RECT 68.02 20.61 69.97 21.01 ;
      RECT 69.31 28.72 69.91 28.92 ;
      RECT 69.71 505.38 69.91 510.01 ;
      RECT 69.31 505.38 69.51 510.01 ;
      RECT 68.71 35.31 69.31 35.51 ;
      RECT 68.79 30.13 69.11 30.73 ;
      RECT 68.79 42.75 69.11 43.35 ;
      RECT 68.91 65.96 69.11 510.01 ;
      RECT 68.07 59.37 68.71 59.97 ;
      RECT 68.51 505.38 68.71 510.01 ;
      RECT 68.11 63.99 68.31 505.18 ;
      RECT 68.11 505.38 68.31 510.01 ;
      RECT 67.51 35.31 68.11 35.51 ;
      RECT 67.86 28.03 68.06 28.77 ;
      RECT 67.71 30.13 68.03 30.73 ;
      RECT 67.71 42.75 68.03 43.35 ;
      RECT 67.71 65.96 67.91 510.01 ;
      RECT 67.61 15.38 67.81 15.98 ;
      RECT 66.81 6.24 67.61 6.84 ;
      RECT 67.31 505.38 67.51 510.01 ;
      RECT 67.11 12.58 67.31 13.85 ;
      RECT 66.91 505.38 67.11 510.01 ;
      RECT 66.31 35.31 66.91 35.51 ;
      RECT 66.61 15.38 66.81 15.98 ;
      RECT 62.95 16.5 66.81 16.7 ;
      RECT 59.53 13.38 66.71 13.58 ;
      RECT 66.39 30.13 66.71 30.73 ;
      RECT 66.39 42.75 66.71 43.35 ;
      RECT 66.36 28.03 66.56 28.77 ;
      RECT 58.41 21.31 66.41 21.51 ;
      RECT 64.45 20.61 66.4 21.01 ;
      RECT 65.71 59.37 66.35 59.97 ;
      RECT 46.21 35.75 66.31 35.95 ;
      RECT 46.21 37.21 66.31 37.41 ;
      RECT 66.11 63.99 66.31 505.18 ;
      RECT 66.11 505.38 66.31 510.01 ;
      RECT 58.66 27.51 66.16 27.71 ;
      RECT 58.66 27.91 66.16 28.11 ;
      RECT 46.21 34.65 66.11 34.85 ;
      RECT 65.71 505.38 65.91 510.01 ;
      RECT 65.11 35.31 65.71 35.51 ;
      RECT 59.13 22.31 65.69 22.51 ;
      RECT 65.31 30.13 65.63 30.73 ;
      RECT 65.31 42.75 65.63 43.35 ;
      RECT 59.33 9.98 65.45 10.18 ;
      RECT 64.37 23.11 65.41 23.31 ;
      RECT 63.91 12.58 65.33 12.78 ;
      RECT 64.31 6.24 65.31 6.84 ;
      RECT 64.51 28.72 65.11 28.92 ;
      RECT 64.91 505.38 65.11 510.01 ;
      RECT 63.13 15.38 64.81 15.58 ;
      RECT 64.21 18.61 64.81 18.81 ;
      RECT 64.51 505.38 64.71 510.01 ;
      RECT 60.25 28.31 64.57 28.51 ;
      RECT 63.91 35.31 64.51 35.51 ;
      RECT 63.99 30.13 64.31 30.73 ;
      RECT 63.99 42.75 64.31 43.35 ;
      RECT 64.11 65.96 64.31 510.01 ;
      RECT 63.95 24.3 64.15 25.07 ;
      RECT 60.75 20.79 64.07 20.99 ;
      RECT 63.27 59.37 63.91 59.97 ;
      RECT 63.71 505.38 63.91 510.01 ;
      RECT 63.21 8.94 63.81 9.14 ;
      RECT 63.31 63.99 63.51 505.18 ;
      RECT 63.31 505.38 63.51 510.01 ;
      RECT 62.71 35.31 63.31 35.51 ;
      RECT 62.91 30.13 63.23 30.73 ;
      RECT 62.91 42.75 63.23 43.35 ;
      RECT 62.91 65.96 63.11 510.01 ;
      RECT 61.29 8.94 63.01 9.14 ;
      RECT 61.85 20.38 62.97 20.58 ;
      RECT 61.41 6.24 62.91 6.84 ;
      RECT 61.81 15.38 62.81 15.72 ;
      RECT 62.51 505.38 62.71 510.01 ;
      RECT 58.01 13.78 62.37 13.98 ;
      RECT 62.11 505.38 62.31 510.01 ;
      RECT 61.51 35.31 62.11 35.51 ;
      RECT 61.59 30.13 61.91 30.73 ;
      RECT 61.59 42.75 61.91 43.35 ;
      RECT 60.91 59.37 61.55 59.97 ;
      RECT 61.31 63.99 61.51 505.18 ;
      RECT 61.31 505.38 61.51 510.01 ;
      RECT 60.14 15.39 61.22 15.59 ;
      RECT 60.91 505.38 61.11 510.01 ;
      RECT 60.41 12.98 61.01 13.18 ;
      RECT 59.01 6.24 60.98 6.84 ;
      RECT 60.31 35.31 60.91 35.51 ;
      RECT 60.67 24.3 60.87 25.07 ;
      RECT 60.51 30.13 60.83 30.73 ;
      RECT 60.51 42.75 60.83 43.35 ;
      RECT 59.85 8.94 60.45 9.14 ;
      RECT 59.41 23.11 60.45 23.31 ;
      RECT 58.42 20.61 60.37 21.01 ;
      RECT 59.71 28.72 60.31 28.92 ;
      RECT 60.11 505.38 60.31 510.01 ;
      RECT 59.71 505.38 59.91 510.01 ;
      RECT 59.11 35.31 59.71 35.51 ;
      RECT 58.66 16.58 59.7 16.78 ;
      RECT 59.19 30.13 59.51 30.73 ;
      RECT 59.19 42.75 59.51 43.35 ;
      RECT 59.31 65.96 59.51 510.01 ;
      RECT 58.47 59.37 59.11 59.97 ;
      RECT 58.91 505.38 59.11 510.01 ;
      RECT 57.91 8.94 58.87 9.14 ;
      RECT 58.51 63.99 58.71 505.18 ;
      RECT 58.51 505.38 58.71 510.01 ;
      RECT 56.61 6.24 58.61 6.84 ;
      RECT 57.91 35.31 58.51 35.51 ;
      RECT 58.26 28.03 58.46 28.77 ;
      RECT 58.11 30.13 58.43 30.73 ;
      RECT 58.11 42.75 58.43 43.35 ;
      RECT 58.11 65.96 58.31 510.01 ;
      RECT 57.71 505.38 57.91 510.01 ;
      RECT 57.17 12.98 57.77 13.18 ;
      RECT 57.31 505.38 57.51 510.01 ;
      RECT 56.71 35.31 57.31 35.51 ;
      RECT 56.79 30.13 57.11 30.73 ;
      RECT 56.79 42.75 57.11 43.35 ;
      RECT 48.71 28.15 56.91 28.75 ;
      RECT 56.11 59.37 56.75 59.97 ;
      RECT 56.51 63.99 56.71 505.18 ;
      RECT 56.51 505.38 56.71 510.01 ;
      RECT 56.11 505.38 56.31 510.01 ;
      RECT 54.21 6.24 56.19 6.84 ;
      RECT 55.51 35.31 56.11 35.51 ;
      RECT 55.71 30.13 56.03 30.73 ;
      RECT 55.71 42.75 56.03 43.35 ;
      RECT 55.31 505.38 55.51 510.01 ;
      RECT 54.91 505.38 55.11 510.01 ;
      RECT 54.31 35.31 54.91 35.51 ;
      RECT 54.39 30.13 54.71 30.73 ;
      RECT 54.39 42.75 54.71 43.35 ;
      RECT 54.51 65.96 54.71 510.01 ;
      RECT 53.67 59.37 54.31 59.97 ;
      RECT 54.11 505.38 54.31 510.01 ;
      RECT 53.71 63.99 53.91 505.18 ;
      RECT 53.71 505.38 53.91 510.01 ;
      RECT 51.81 6.24 53.79 6.84 ;
      RECT 53.11 35.31 53.71 35.51 ;
      RECT 53.31 30.13 53.63 30.73 ;
      RECT 53.31 42.75 53.63 43.35 ;
      RECT 52.11 15.51 53.51 15.71 ;
      RECT 53.31 65.96 53.51 510.01 ;
      RECT 52.91 505.38 53.11 510.01 ;
      RECT 52.51 505.38 52.71 510.01 ;
      RECT 51.91 35.31 52.51 35.51 ;
      RECT 51.99 30.13 52.31 30.73 ;
      RECT 51.99 42.75 52.31 43.35 ;
      RECT 51.31 59.37 51.95 59.97 ;
      RECT 51.71 63.99 51.91 505.18 ;
      RECT 51.71 505.38 51.91 510.01 ;
      RECT 51.31 505.38 51.51 510.01 ;
      RECT 49.41 6.24 51.39 6.84 ;
      RECT 50.71 35.31 51.31 35.51 ;
      RECT 50.91 30.13 51.23 30.73 ;
      RECT 50.91 42.75 51.23 43.35 ;
      RECT 50.51 505.38 50.71 510.01 ;
      RECT 50.11 505.38 50.31 510.01 ;
      RECT 49.51 35.31 50.11 35.51 ;
      RECT 49.59 30.13 49.91 30.73 ;
      RECT 49.59 42.75 49.91 43.35 ;
      RECT 49.71 65.96 49.91 510.01 ;
      RECT 48.87 59.37 49.51 59.97 ;
      RECT 49.31 505.38 49.51 510.01 ;
      RECT 48.91 63.99 49.11 505.18 ;
      RECT 48.91 505.38 49.11 510.01 ;
      RECT 47.61 6.24 49.01 6.84 ;
      RECT 48.31 35.31 48.91 35.51 ;
      RECT 48.51 30.13 48.83 30.73 ;
      RECT 48.51 42.75 48.83 43.35 ;
      RECT 48.51 65.96 48.71 510.01 ;
      RECT 48.11 505.38 48.31 510.01 ;
      RECT 47.31 68.76 47.51 70.14 ;
      RECT 47.31 70.34 47.51 71.16 ;
      RECT 47.31 71.36 47.51 72.18 ;
      RECT 47.31 72.38 47.51 73.54 ;
      RECT 47.31 73.74 47.51 74.56 ;
      RECT 47.31 74.76 47.51 75.58 ;
      RECT 47.31 75.78 47.51 76.94 ;
      RECT 47.31 77.14 47.51 77.96 ;
      RECT 47.31 78.16 47.51 78.98 ;
      RECT 47.31 79.18 47.51 80.34 ;
      RECT 47.31 80.54 47.51 81.36 ;
      RECT 47.31 81.56 47.51 82.38 ;
      RECT 47.31 82.58 47.51 83.74 ;
      RECT 47.31 83.94 47.51 84.76 ;
      RECT 47.31 84.96 47.51 85.78 ;
      RECT 47.31 85.98 47.51 87.14 ;
      RECT 47.31 87.34 47.51 88.16 ;
      RECT 47.31 88.36 47.51 89.18 ;
      RECT 47.31 89.38 47.51 90.54 ;
      RECT 47.31 90.74 47.51 91.56 ;
      RECT 47.31 91.76 47.51 92.58 ;
      RECT 47.31 92.78 47.51 93.94 ;
      RECT 47.31 94.14 47.51 94.96 ;
      RECT 47.31 95.16 47.51 95.98 ;
      RECT 47.31 96.18 47.51 97.34 ;
      RECT 47.31 97.54 47.51 98.36 ;
      RECT 47.31 98.56 47.51 99.38 ;
      RECT 47.31 99.58 47.51 100.74 ;
      RECT 47.31 100.94 47.51 101.76 ;
      RECT 47.31 101.96 47.51 102.78 ;
      RECT 47.31 102.98 47.51 104.14 ;
      RECT 47.31 104.34 47.51 105.16 ;
      RECT 47.31 105.36 47.51 106.18 ;
      RECT 47.31 106.38 47.51 107.54 ;
      RECT 47.31 107.74 47.51 108.56 ;
      RECT 47.31 108.76 47.51 109.58 ;
      RECT 47.31 109.78 47.51 110.94 ;
      RECT 47.31 111.14 47.51 111.96 ;
      RECT 47.31 112.16 47.51 112.98 ;
      RECT 47.31 113.18 47.51 114.34 ;
      RECT 47.31 114.54 47.51 115.36 ;
      RECT 47.31 115.56 47.51 116.38 ;
      RECT 47.31 116.58 47.51 117.74 ;
      RECT 47.31 117.94 47.51 118.76 ;
      RECT 47.31 118.96 47.51 119.78 ;
      RECT 47.31 119.98 47.51 121.14 ;
      RECT 47.31 121.34 47.51 122.16 ;
      RECT 47.31 122.36 47.51 123.18 ;
      RECT 47.31 123.38 47.51 124.54 ;
      RECT 47.31 124.74 47.51 125.56 ;
      RECT 47.31 125.76 47.51 126.58 ;
      RECT 47.31 126.78 47.51 127.94 ;
      RECT 47.31 128.14 47.51 128.96 ;
      RECT 47.31 129.16 47.51 129.98 ;
      RECT 47.31 130.18 47.51 131.34 ;
      RECT 47.31 131.54 47.51 132.36 ;
      RECT 47.31 132.56 47.51 133.38 ;
      RECT 47.31 133.58 47.51 134.74 ;
      RECT 47.31 134.94 47.51 135.76 ;
      RECT 47.31 135.96 47.51 136.78 ;
      RECT 47.31 136.98 47.51 138.14 ;
      RECT 47.31 138.34 47.51 139.16 ;
      RECT 47.31 139.36 47.51 140.18 ;
      RECT 47.31 140.38 47.51 141.54 ;
      RECT 47.31 141.74 47.51 142.56 ;
      RECT 47.31 142.76 47.51 143.58 ;
      RECT 47.31 143.78 47.51 144.94 ;
      RECT 47.31 145.14 47.51 145.96 ;
      RECT 47.31 146.16 47.51 146.98 ;
      RECT 47.31 147.18 47.51 148.34 ;
      RECT 47.31 148.54 47.51 149.36 ;
      RECT 47.31 149.56 47.51 150.38 ;
      RECT 47.31 150.58 47.51 151.74 ;
      RECT 47.31 151.94 47.51 152.76 ;
      RECT 47.31 152.96 47.51 153.78 ;
      RECT 47.31 153.98 47.51 155.14 ;
      RECT 47.31 155.34 47.51 156.16 ;
      RECT 47.31 156.36 47.51 157.18 ;
      RECT 47.31 157.38 47.51 158.54 ;
      RECT 47.31 158.74 47.51 159.56 ;
      RECT 47.31 159.76 47.51 160.58 ;
      RECT 47.31 160.78 47.51 161.94 ;
      RECT 47.31 162.14 47.51 162.96 ;
      RECT 47.31 163.16 47.51 163.98 ;
      RECT 47.31 164.18 47.51 165.34 ;
      RECT 47.31 165.54 47.51 166.36 ;
      RECT 47.31 166.56 47.51 167.38 ;
      RECT 47.31 167.58 47.51 168.74 ;
      RECT 47.31 168.94 47.51 169.76 ;
      RECT 47.31 169.96 47.51 170.78 ;
      RECT 47.31 170.98 47.51 172.14 ;
      RECT 47.31 172.34 47.51 173.16 ;
      RECT 47.31 173.36 47.51 174.18 ;
      RECT 47.31 174.38 47.51 175.54 ;
      RECT 47.31 175.74 47.51 176.56 ;
      RECT 47.31 176.76 47.51 177.58 ;
      RECT 47.31 177.78 47.51 178.94 ;
      RECT 47.31 179.14 47.51 179.96 ;
      RECT 47.31 180.16 47.51 180.98 ;
      RECT 47.31 181.18 47.51 182.34 ;
      RECT 47.31 182.54 47.51 183.36 ;
      RECT 47.31 183.56 47.51 184.38 ;
      RECT 47.31 184.58 47.51 185.74 ;
      RECT 47.31 185.94 47.51 186.76 ;
      RECT 47.31 186.96 47.51 187.78 ;
      RECT 47.31 187.98 47.51 189.14 ;
      RECT 47.31 189.34 47.51 190.16 ;
      RECT 47.31 190.36 47.51 191.18 ;
      RECT 47.31 191.38 47.51 192.54 ;
      RECT 47.31 192.74 47.51 193.56 ;
      RECT 47.31 193.76 47.51 194.58 ;
      RECT 47.31 194.78 47.51 195.94 ;
      RECT 47.31 196.14 47.51 196.96 ;
      RECT 47.31 197.16 47.51 197.98 ;
      RECT 47.31 198.18 47.51 199.34 ;
      RECT 47.31 199.54 47.51 200.36 ;
      RECT 47.31 200.56 47.51 201.38 ;
      RECT 47.31 201.58 47.51 202.74 ;
      RECT 47.31 202.94 47.51 203.76 ;
      RECT 47.31 203.96 47.51 204.78 ;
      RECT 47.31 204.98 47.51 206.14 ;
      RECT 47.31 206.34 47.51 207.16 ;
      RECT 47.31 207.36 47.51 208.18 ;
      RECT 47.31 208.38 47.51 209.54 ;
      RECT 47.31 209.74 47.51 210.56 ;
      RECT 47.31 210.76 47.51 211.58 ;
      RECT 47.31 211.78 47.51 212.94 ;
      RECT 47.31 213.14 47.51 213.96 ;
      RECT 47.31 214.16 47.51 214.98 ;
      RECT 47.31 215.18 47.51 216.34 ;
      RECT 47.31 216.54 47.51 217.36 ;
      RECT 47.31 217.56 47.51 218.38 ;
      RECT 47.31 218.58 47.51 219.74 ;
      RECT 47.31 219.94 47.51 220.76 ;
      RECT 47.31 220.96 47.51 221.78 ;
      RECT 47.31 221.98 47.51 223.14 ;
      RECT 47.31 223.34 47.51 224.16 ;
      RECT 47.31 224.36 47.51 225.18 ;
      RECT 47.31 225.38 47.51 226.54 ;
      RECT 47.31 226.74 47.51 227.56 ;
      RECT 47.31 227.76 47.51 228.58 ;
      RECT 47.31 228.78 47.51 229.94 ;
      RECT 47.31 230.14 47.51 230.96 ;
      RECT 47.31 231.16 47.51 231.98 ;
      RECT 47.31 232.18 47.51 233.34 ;
      RECT 47.31 233.54 47.51 234.36 ;
      RECT 47.31 234.56 47.51 235.38 ;
      RECT 47.31 235.58 47.51 236.74 ;
      RECT 47.31 236.94 47.51 237.76 ;
      RECT 47.31 237.96 47.51 238.78 ;
      RECT 47.31 238.98 47.51 240.14 ;
      RECT 47.31 240.34 47.51 241.16 ;
      RECT 47.31 241.36 47.51 242.18 ;
      RECT 47.31 242.38 47.51 243.54 ;
      RECT 47.31 243.74 47.51 244.56 ;
      RECT 47.31 244.76 47.51 245.58 ;
      RECT 47.31 245.78 47.51 246.94 ;
      RECT 47.31 247.14 47.51 247.96 ;
      RECT 47.31 248.16 47.51 248.98 ;
      RECT 47.31 249.18 47.51 250.34 ;
      RECT 47.31 250.54 47.51 251.36 ;
      RECT 47.31 251.56 47.51 252.38 ;
      RECT 47.31 252.58 47.51 253.74 ;
      RECT 47.31 253.94 47.51 254.76 ;
      RECT 47.31 254.96 47.51 255.78 ;
      RECT 47.31 255.98 47.51 257.14 ;
      RECT 47.31 257.34 47.51 258.16 ;
      RECT 47.31 258.36 47.51 259.18 ;
      RECT 47.31 259.38 47.51 260.54 ;
      RECT 47.31 260.74 47.51 261.56 ;
      RECT 47.31 261.76 47.51 262.58 ;
      RECT 47.31 262.78 47.51 263.94 ;
      RECT 47.31 264.14 47.51 264.96 ;
      RECT 47.31 265.16 47.51 265.98 ;
      RECT 47.31 266.18 47.51 267.34 ;
      RECT 47.31 267.54 47.51 268.36 ;
      RECT 47.31 268.56 47.51 269.38 ;
      RECT 47.31 269.58 47.51 270.74 ;
      RECT 47.31 270.94 47.51 271.76 ;
      RECT 47.31 271.96 47.51 272.78 ;
      RECT 47.31 272.98 47.51 274.14 ;
      RECT 47.31 274.34 47.51 275.16 ;
      RECT 47.31 275.36 47.51 276.18 ;
      RECT 47.31 276.38 47.51 277.54 ;
      RECT 47.31 277.74 47.51 278.56 ;
      RECT 47.31 278.76 47.51 279.58 ;
      RECT 47.31 279.78 47.51 280.94 ;
      RECT 47.31 281.14 47.51 281.96 ;
      RECT 47.31 282.16 47.51 282.98 ;
      RECT 47.31 283.18 47.51 284.34 ;
      RECT 47.31 284.54 47.51 285.36 ;
      RECT 47.31 285.56 47.51 286.38 ;
      RECT 47.31 286.58 47.51 287.74 ;
      RECT 47.31 287.94 47.51 288.76 ;
      RECT 47.31 288.96 47.51 289.78 ;
      RECT 47.31 289.98 47.51 291.14 ;
      RECT 47.31 291.34 47.51 292.16 ;
      RECT 47.31 292.36 47.51 293.18 ;
      RECT 47.31 293.38 47.51 294.54 ;
      RECT 47.31 294.74 47.51 295.56 ;
      RECT 47.31 295.76 47.51 296.58 ;
      RECT 47.31 296.78 47.51 297.94 ;
      RECT 47.31 298.14 47.51 298.96 ;
      RECT 47.31 299.16 47.51 299.98 ;
      RECT 47.31 300.18 47.51 301.34 ;
      RECT 47.31 301.54 47.51 302.36 ;
      RECT 47.31 302.56 47.51 303.38 ;
      RECT 47.31 303.58 47.51 304.74 ;
      RECT 47.31 304.94 47.51 305.76 ;
      RECT 47.31 305.96 47.51 306.78 ;
      RECT 47.31 306.98 47.51 308.14 ;
      RECT 47.31 308.34 47.51 309.16 ;
      RECT 47.31 309.36 47.51 310.18 ;
      RECT 47.31 310.38 47.51 311.54 ;
      RECT 47.31 311.74 47.51 312.56 ;
      RECT 47.31 312.76 47.51 313.58 ;
      RECT 47.31 313.78 47.51 314.94 ;
      RECT 47.31 315.14 47.51 315.96 ;
      RECT 47.31 316.16 47.51 316.98 ;
      RECT 47.31 317.18 47.51 318.34 ;
      RECT 47.31 318.54 47.51 319.36 ;
      RECT 47.31 319.56 47.51 320.38 ;
      RECT 47.31 320.58 47.51 321.74 ;
      RECT 47.31 321.94 47.51 322.76 ;
      RECT 47.31 322.96 47.51 323.78 ;
      RECT 47.31 323.98 47.51 325.14 ;
      RECT 47.31 325.34 47.51 326.16 ;
      RECT 47.31 326.36 47.51 327.18 ;
      RECT 47.31 327.38 47.51 328.54 ;
      RECT 47.31 328.74 47.51 329.56 ;
      RECT 47.31 329.76 47.51 330.58 ;
      RECT 47.31 330.78 47.51 331.94 ;
      RECT 47.31 332.14 47.51 332.96 ;
      RECT 47.31 333.16 47.51 333.98 ;
      RECT 47.31 334.18 47.51 335.34 ;
      RECT 47.31 335.54 47.51 336.36 ;
      RECT 47.31 336.56 47.51 337.38 ;
      RECT 47.31 337.58 47.51 338.74 ;
      RECT 47.31 338.94 47.51 339.76 ;
      RECT 47.31 339.96 47.51 340.78 ;
      RECT 47.31 340.98 47.51 342.14 ;
      RECT 47.31 342.34 47.51 343.16 ;
      RECT 47.31 343.36 47.51 344.18 ;
      RECT 47.31 344.38 47.51 345.54 ;
      RECT 47.31 345.74 47.51 346.56 ;
      RECT 47.31 346.76 47.51 347.58 ;
      RECT 47.31 347.78 47.51 348.94 ;
      RECT 47.31 349.14 47.51 349.96 ;
      RECT 47.31 350.16 47.51 350.98 ;
      RECT 47.31 351.18 47.51 352.34 ;
      RECT 47.31 352.54 47.51 353.36 ;
      RECT 47.31 353.56 47.51 354.38 ;
      RECT 47.31 354.58 47.51 355.74 ;
      RECT 47.31 355.94 47.51 356.76 ;
      RECT 47.31 356.96 47.51 357.78 ;
      RECT 47.31 357.98 47.51 359.14 ;
      RECT 47.31 359.34 47.51 360.16 ;
      RECT 47.31 360.36 47.51 361.18 ;
      RECT 47.31 361.38 47.51 362.54 ;
      RECT 47.31 362.74 47.51 363.56 ;
      RECT 47.31 363.76 47.51 364.58 ;
      RECT 47.31 364.78 47.51 365.94 ;
      RECT 47.31 366.14 47.51 366.96 ;
      RECT 47.31 367.16 47.51 367.98 ;
      RECT 47.31 368.18 47.51 369.34 ;
      RECT 47.31 369.54 47.51 370.36 ;
      RECT 47.31 370.56 47.51 371.38 ;
      RECT 47.31 371.58 47.51 372.74 ;
      RECT 47.31 372.94 47.51 373.76 ;
      RECT 47.31 373.96 47.51 374.78 ;
      RECT 47.31 374.98 47.51 376.14 ;
      RECT 47.31 376.34 47.51 377.16 ;
      RECT 47.31 377.36 47.51 378.18 ;
      RECT 47.31 378.38 47.51 379.54 ;
      RECT 47.31 379.74 47.51 380.56 ;
      RECT 47.31 380.76 47.51 381.58 ;
      RECT 47.31 381.78 47.51 382.94 ;
      RECT 47.31 383.14 47.51 383.96 ;
      RECT 47.31 384.16 47.51 384.98 ;
      RECT 47.31 385.18 47.51 386.34 ;
      RECT 47.31 386.54 47.51 387.36 ;
      RECT 47.31 387.56 47.51 388.38 ;
      RECT 47.31 388.58 47.51 389.74 ;
      RECT 47.31 389.94 47.51 390.76 ;
      RECT 47.31 390.96 47.51 391.78 ;
      RECT 47.31 391.98 47.51 393.14 ;
      RECT 47.31 393.34 47.51 394.16 ;
      RECT 47.31 394.36 47.51 395.18 ;
      RECT 47.31 395.38 47.51 396.54 ;
      RECT 47.31 396.74 47.51 397.56 ;
      RECT 47.31 397.76 47.51 398.58 ;
      RECT 47.31 398.78 47.51 399.94 ;
      RECT 47.31 400.14 47.51 400.96 ;
      RECT 47.31 401.16 47.51 401.98 ;
      RECT 47.31 402.18 47.51 403.34 ;
      RECT 47.31 403.54 47.51 404.36 ;
      RECT 47.31 404.56 47.51 405.38 ;
      RECT 47.31 405.58 47.51 406.74 ;
      RECT 47.31 406.94 47.51 407.76 ;
      RECT 47.31 407.96 47.51 408.78 ;
      RECT 47.31 408.98 47.51 410.14 ;
      RECT 47.31 410.34 47.51 411.16 ;
      RECT 47.31 411.36 47.51 412.18 ;
      RECT 47.31 412.38 47.51 413.54 ;
      RECT 47.31 413.74 47.51 414.56 ;
      RECT 47.31 414.76 47.51 415.58 ;
      RECT 47.31 415.78 47.51 416.94 ;
      RECT 47.31 417.14 47.51 417.96 ;
      RECT 47.31 418.16 47.51 418.98 ;
      RECT 47.31 419.18 47.51 420.34 ;
      RECT 47.31 420.54 47.51 421.36 ;
      RECT 47.31 421.56 47.51 422.38 ;
      RECT 47.31 422.58 47.51 423.74 ;
      RECT 47.31 423.94 47.51 424.76 ;
      RECT 47.31 424.96 47.51 425.78 ;
      RECT 47.31 425.98 47.51 427.14 ;
      RECT 47.31 427.34 47.51 428.16 ;
      RECT 47.31 428.36 47.51 429.18 ;
      RECT 47.31 429.38 47.51 430.54 ;
      RECT 47.31 430.74 47.51 431.56 ;
      RECT 47.31 431.76 47.51 432.58 ;
      RECT 47.31 432.78 47.51 433.94 ;
      RECT 47.31 434.14 47.51 434.96 ;
      RECT 47.31 435.16 47.51 435.98 ;
      RECT 47.31 436.18 47.51 437.34 ;
      RECT 47.31 437.54 47.51 438.36 ;
      RECT 47.31 438.56 47.51 439.38 ;
      RECT 47.31 439.58 47.51 440.74 ;
      RECT 47.31 440.94 47.51 441.76 ;
      RECT 47.31 441.96 47.51 442.78 ;
      RECT 47.31 442.98 47.51 444.14 ;
      RECT 47.31 444.34 47.51 445.16 ;
      RECT 47.31 445.36 47.51 446.18 ;
      RECT 47.31 446.38 47.51 447.54 ;
      RECT 47.31 447.74 47.51 448.56 ;
      RECT 47.31 448.76 47.51 449.58 ;
      RECT 47.31 449.78 47.51 450.94 ;
      RECT 47.31 451.14 47.51 451.96 ;
      RECT 47.31 452.16 47.51 452.98 ;
      RECT 47.31 453.18 47.51 454.34 ;
      RECT 47.31 454.54 47.51 455.36 ;
      RECT 47.31 455.56 47.51 456.38 ;
      RECT 47.31 456.58 47.51 457.74 ;
      RECT 47.31 457.94 47.51 458.76 ;
      RECT 47.31 458.96 47.51 459.78 ;
      RECT 47.31 459.98 47.51 461.14 ;
      RECT 47.31 461.34 47.51 462.16 ;
      RECT 47.31 462.36 47.51 463.18 ;
      RECT 47.31 463.38 47.51 464.54 ;
      RECT 47.31 464.74 47.51 465.56 ;
      RECT 47.31 465.76 47.51 466.58 ;
      RECT 47.31 466.78 47.51 467.94 ;
      RECT 47.31 468.14 47.51 468.96 ;
      RECT 47.31 469.16 47.51 469.98 ;
      RECT 47.31 470.18 47.51 471.34 ;
      RECT 47.31 471.54 47.51 472.36 ;
      RECT 47.31 472.56 47.51 473.38 ;
      RECT 47.31 473.58 47.51 474.74 ;
      RECT 47.31 474.94 47.51 475.76 ;
      RECT 47.31 475.96 47.51 476.78 ;
      RECT 47.31 476.98 47.51 478.14 ;
      RECT 47.31 478.34 47.51 479.16 ;
      RECT 47.31 479.36 47.51 480.18 ;
      RECT 47.31 480.38 47.51 481.54 ;
      RECT 47.31 481.74 47.51 482.56 ;
      RECT 47.31 482.76 47.51 483.58 ;
      RECT 47.31 483.78 47.51 484.94 ;
      RECT 47.31 485.14 47.51 485.96 ;
      RECT 47.31 486.16 47.51 486.98 ;
      RECT 47.31 487.18 47.51 488.34 ;
      RECT 47.31 488.54 47.51 489.36 ;
      RECT 47.31 489.56 47.51 490.38 ;
      RECT 47.31 490.58 47.51 491.74 ;
      RECT 47.31 491.94 47.51 492.76 ;
      RECT 47.31 492.96 47.51 493.78 ;
      RECT 47.31 493.98 47.51 495.14 ;
      RECT 47.31 495.34 47.51 496.16 ;
      RECT 47.31 496.36 47.51 497.18 ;
      RECT 47.31 497.38 47.51 498.54 ;
      RECT 47.31 498.74 47.51 499.56 ;
      RECT 47.31 499.76 47.51 500.58 ;
      RECT 47.31 500.78 47.51 501.94 ;
      RECT 47.31 502.14 47.51 502.96 ;
      RECT 47.31 503.16 47.51 503.98 ;
      RECT 47.31 504.18 47.51 506.38 ;
      RECT 47.31 506.58 47.51 507.4 ;
      RECT 47.31 507.6 47.51 508.42 ;
      RECT 47.31 508.62 47.51 510 ;
      RECT 45.81 6.24 47.21 6.84 ;
      RECT 46.51 505.38 46.71 510.01 ;
      RECT 45.91 35.31 46.51 35.51 ;
      RECT 45.99 30.13 46.31 30.73 ;
      RECT 45.99 42.75 46.31 43.35 ;
      RECT 37.91 28.15 46.11 28.75 ;
      RECT 45.31 59.37 45.95 59.97 ;
      RECT 27.01 35.75 45.91 35.95 ;
      RECT 27.01 37.21 45.91 37.41 ;
      RECT 45.71 63.99 45.91 505.18 ;
      RECT 45.71 505.38 45.91 510.01 ;
      RECT 27.01 34.65 45.71 34.85 ;
      RECT 45.31 505.38 45.51 510.01 ;
      RECT 43.43 6.24 45.41 6.84 ;
      RECT 44.71 35.31 45.31 35.51 ;
      RECT 44.91 30.13 45.23 30.73 ;
      RECT 44.91 42.75 45.23 43.35 ;
      RECT 44.51 505.38 44.71 510.01 ;
      RECT 44.11 505.38 44.31 510.01 ;
      RECT 43.51 35.31 44.11 35.51 ;
      RECT 43.59 30.13 43.91 30.73 ;
      RECT 43.59 42.75 43.91 43.35 ;
      RECT 43.71 65.96 43.91 510.01 ;
      RECT 42.87 59.37 43.51 59.97 ;
      RECT 43.31 505.38 43.51 510.01 ;
      RECT 42.91 63.99 43.11 505.18 ;
      RECT 42.91 505.38 43.11 510.01 ;
      RECT 41.03 6.24 43.01 6.84 ;
      RECT 42.31 35.31 42.91 35.51 ;
      RECT 42.51 30.13 42.83 30.73 ;
      RECT 42.51 42.75 42.83 43.35 ;
      RECT 41.31 15.51 42.71 15.71 ;
      RECT 42.51 65.96 42.71 510.01 ;
      RECT 42.11 505.38 42.31 510.01 ;
      RECT 41.71 505.38 41.91 510.01 ;
      RECT 41.11 35.31 41.71 35.51 ;
      RECT 41.19 30.13 41.51 30.73 ;
      RECT 41.19 42.75 41.51 43.35 ;
      RECT 40.51 59.37 41.15 59.97 ;
      RECT 40.91 63.99 41.11 505.18 ;
      RECT 40.91 505.38 41.11 510.01 ;
      RECT 40.51 505.38 40.71 510.01 ;
      RECT 38.63 6.24 40.61 6.84 ;
      RECT 39.91 35.31 40.51 35.51 ;
      RECT 40.11 30.13 40.43 30.73 ;
      RECT 40.11 42.75 40.43 43.35 ;
      RECT 39.71 505.38 39.91 510.01 ;
      RECT 39.31 505.38 39.51 510.01 ;
      RECT 38.71 35.31 39.31 35.51 ;
      RECT 38.79 30.13 39.11 30.73 ;
      RECT 38.79 42.75 39.11 43.35 ;
      RECT 38.91 65.96 39.11 510.01 ;
      RECT 38.07 59.37 38.71 59.97 ;
      RECT 38.51 505.38 38.71 510.01 ;
      RECT 38.11 63.99 38.31 505.18 ;
      RECT 38.11 505.38 38.31 510.01 ;
      RECT 36.21 6.24 38.21 6.84 ;
      RECT 37.51 35.31 38.11 35.51 ;
      RECT 37.71 30.13 38.03 30.73 ;
      RECT 37.71 42.75 38.03 43.35 ;
      RECT 37.71 65.96 37.91 510.01 ;
      RECT 37.05 12.98 37.65 13.18 ;
      RECT 37.31 505.38 37.51 510.01 ;
      RECT 36.91 505.38 37.11 510.01 ;
      RECT 35.95 8.94 36.91 9.14 ;
      RECT 36.31 35.31 36.91 35.51 ;
      RECT 32.45 13.78 36.81 13.98 ;
      RECT 36.39 30.13 36.71 30.73 ;
      RECT 36.39 42.75 36.71 43.35 ;
      RECT 36.36 28.03 36.56 28.77 ;
      RECT 28.41 21.31 36.41 21.51 ;
      RECT 34.45 20.61 36.4 21.01 ;
      RECT 35.71 59.37 36.35 59.97 ;
      RECT 36.11 63.99 36.31 505.18 ;
      RECT 36.11 505.38 36.31 510.01 ;
      RECT 35.12 16.58 36.16 16.78 ;
      RECT 28.66 27.51 36.16 27.71 ;
      RECT 28.66 27.91 36.16 28.11 ;
      RECT 35.71 505.38 35.91 510.01 ;
      RECT 33.84 6.24 35.81 6.84 ;
      RECT 35.11 35.31 35.71 35.51 ;
      RECT 29.13 22.31 35.69 22.51 ;
      RECT 35.31 30.13 35.63 30.73 ;
      RECT 35.31 42.75 35.63 43.35 ;
      RECT 29.37 9.98 35.49 10.18 ;
      RECT 34.37 23.11 35.41 23.31 ;
      RECT 28.11 13.38 35.29 13.58 ;
      RECT 34.51 28.72 35.11 28.92 ;
      RECT 34.91 505.38 35.11 510.01 ;
      RECT 34.37 8.94 34.97 9.14 ;
      RECT 34.51 505.38 34.71 510.01 ;
      RECT 33.6 15.39 34.68 15.59 ;
      RECT 30.25 28.31 34.57 28.51 ;
      RECT 33.91 35.31 34.51 35.51 ;
      RECT 33.81 12.98 34.41 13.18 ;
      RECT 33.99 30.13 34.31 30.73 ;
      RECT 33.99 42.75 34.31 43.35 ;
      RECT 34.11 65.96 34.31 510.01 ;
      RECT 33.95 24.3 34.15 25.07 ;
      RECT 30.75 20.79 34.07 20.99 ;
      RECT 33.27 59.37 33.91 59.97 ;
      RECT 33.71 505.38 33.91 510.01 ;
      RECT 31.81 8.94 33.53 9.14 ;
      RECT 33.31 63.99 33.51 505.18 ;
      RECT 33.31 505.38 33.51 510.01 ;
      RECT 31.91 6.24 33.41 6.84 ;
      RECT 32.71 35.31 33.31 35.51 ;
      RECT 32.91 30.13 33.23 30.73 ;
      RECT 32.91 42.75 33.23 43.35 ;
      RECT 32.91 65.96 33.11 510.01 ;
      RECT 32.01 15.38 33.01 15.72 ;
      RECT 31.85 20.38 32.97 20.58 ;
      RECT 32.51 505.38 32.71 510.01 ;
      RECT 32.11 505.38 32.31 510.01 ;
      RECT 31.51 35.31 32.11 35.51 ;
      RECT 31.59 30.13 31.91 30.73 ;
      RECT 31.59 42.75 31.91 43.35 ;
      RECT 28.01 16.5 31.87 16.7 ;
      RECT 30.01 15.38 31.69 15.58 ;
      RECT 31.01 8.94 31.61 9.14 ;
      RECT 30.91 59.37 31.55 59.97 ;
      RECT 31.31 63.99 31.51 505.18 ;
      RECT 31.31 505.38 31.51 510.01 ;
      RECT 30.91 505.38 31.11 510.01 ;
      RECT 29.49 12.58 30.91 12.78 ;
      RECT 30.31 35.31 30.91 35.51 ;
      RECT 30.67 24.3 30.87 25.07 ;
      RECT 30.51 30.13 30.83 30.73 ;
      RECT 30.51 42.75 30.83 43.35 ;
      RECT 30.01 18.61 30.61 18.81 ;
      RECT 29.51 6.24 30.51 6.84 ;
      RECT 29.41 23.11 30.45 23.31 ;
      RECT 28.42 20.61 30.37 21.01 ;
      RECT 29.71 28.72 30.31 28.92 ;
      RECT 30.11 505.38 30.31 510.01 ;
      RECT 29.71 505.38 29.91 510.01 ;
      RECT 29.11 35.31 29.71 35.51 ;
      RECT 29.19 30.13 29.51 30.73 ;
      RECT 29.19 42.75 29.51 43.35 ;
      RECT 29.31 65.96 29.51 510.01 ;
      RECT 28.47 59.37 29.11 59.97 ;
      RECT 28.91 505.38 29.11 510.01 ;
      RECT 28.51 63.99 28.71 505.18 ;
      RECT 28.51 505.38 28.71 510.01 ;
      RECT 27.91 35.31 28.51 35.51 ;
      RECT 28.26 28.03 28.46 28.77 ;
      RECT 28.11 30.13 28.43 30.73 ;
      RECT 28.11 42.75 28.43 43.35 ;
      RECT 28.11 65.96 28.31 510.01 ;
      RECT 28.01 15.38 28.21 15.98 ;
      RECT 27.21 6.24 28.01 6.84 ;
      RECT 27.71 505.38 27.91 510.01 ;
      RECT 27.51 12.58 27.71 13.85 ;
      RECT 27.31 505.38 27.51 510.01 ;
      RECT 26.71 35.31 27.31 35.51 ;
      RECT 27.01 15.38 27.21 15.98 ;
      RECT 23.35 16.5 27.21 16.7 ;
      RECT 19.93 13.38 27.11 13.58 ;
      RECT 26.79 30.13 27.11 30.73 ;
      RECT 26.79 42.75 27.11 43.35 ;
      RECT 26.76 28.03 26.96 28.77 ;
      RECT 18.81 21.31 26.81 21.51 ;
      RECT 24.85 20.61 26.8 21.01 ;
      RECT 26.11 59.37 26.75 59.97 ;
      RECT 7.81 35.75 26.71 35.95 ;
      RECT 7.81 37.21 26.71 37.41 ;
      RECT 26.51 63.99 26.71 505.18 ;
      RECT 26.51 505.38 26.71 510.01 ;
      RECT 19.06 27.51 26.56 27.71 ;
      RECT 19.06 27.91 26.56 28.11 ;
      RECT 7.81 34.65 26.51 34.85 ;
      RECT 26.11 505.38 26.31 510.01 ;
      RECT 25.51 35.31 26.11 35.51 ;
      RECT 19.53 22.31 26.09 22.51 ;
      RECT 25.71 30.13 26.03 30.73 ;
      RECT 25.71 42.75 26.03 43.35 ;
      RECT 19.73 9.98 25.85 10.18 ;
      RECT 24.77 23.11 25.81 23.31 ;
      RECT 24.31 12.58 25.73 12.78 ;
      RECT 24.71 6.24 25.71 6.84 ;
      RECT 24.91 28.72 25.51 28.92 ;
      RECT 25.31 505.38 25.51 510.01 ;
      RECT 23.53 15.38 25.21 15.58 ;
      RECT 24.61 18.61 25.21 18.81 ;
      RECT 24.91 505.38 25.11 510.01 ;
      RECT 20.65 28.31 24.97 28.51 ;
      RECT 24.31 35.31 24.91 35.51 ;
      RECT 24.39 30.13 24.71 30.73 ;
      RECT 24.39 42.75 24.71 43.35 ;
      RECT 24.51 65.96 24.71 510.01 ;
      RECT 24.35 24.3 24.55 25.07 ;
      RECT 21.15 20.79 24.47 20.99 ;
      RECT 23.67 59.37 24.31 59.97 ;
      RECT 24.11 505.38 24.31 510.01 ;
      RECT 23.61 8.94 24.21 9.14 ;
      RECT 23.71 63.99 23.91 505.18 ;
      RECT 23.71 505.38 23.91 510.01 ;
      RECT 23.11 35.31 23.71 35.51 ;
      RECT 23.31 30.13 23.63 30.73 ;
      RECT 23.31 42.75 23.63 43.35 ;
      RECT 23.31 65.96 23.51 510.01 ;
      RECT 21.69 8.94 23.41 9.14 ;
      RECT 22.25 20.38 23.37 20.58 ;
      RECT 21.81 6.24 23.31 6.84 ;
      RECT 22.21 15.38 23.21 15.72 ;
      RECT 22.91 505.38 23.11 510.01 ;
      RECT 18.41 13.78 22.77 13.98 ;
      RECT 22.51 505.38 22.71 510.01 ;
      RECT 21.91 35.31 22.51 35.51 ;
      RECT 21.99 30.13 22.31 30.73 ;
      RECT 21.99 42.75 22.31 43.35 ;
      RECT 21.31 59.37 21.95 59.97 ;
      RECT 21.71 63.99 21.91 505.18 ;
      RECT 21.71 505.38 21.91 510.01 ;
      RECT 20.54 15.39 21.62 15.59 ;
      RECT 21.31 505.38 21.51 510.01 ;
      RECT 19.81 6.24 21.41 6.84 ;
      RECT 20.81 12.98 21.41 13.18 ;
      RECT 20.71 35.31 21.31 35.51 ;
      RECT 21.07 24.3 21.27 25.07 ;
      RECT 20.91 30.13 21.23 30.73 ;
      RECT 20.91 42.75 21.23 43.35 ;
      RECT 20.25 8.94 20.85 9.14 ;
      RECT 19.81 23.11 20.85 23.31 ;
      RECT 18.82 20.61 20.77 21.01 ;
      RECT 20.11 28.72 20.71 28.92 ;
      RECT 20.51 505.38 20.71 510.01 ;
      RECT 20.11 505.38 20.31 510.01 ;
      RECT 19.51 35.31 20.11 35.51 ;
      RECT 19.06 16.58 20.1 16.78 ;
      RECT 19.59 30.13 19.91 30.73 ;
      RECT 19.59 42.75 19.91 43.35 ;
      RECT 19.71 65.96 19.91 510.01 ;
      RECT 18.87 59.37 19.51 59.97 ;
      RECT 19.31 505.38 19.51 510.01 ;
      RECT 18.81 6.24 19.41 6.84 ;
      RECT 18.31 8.94 19.27 9.14 ;
      RECT 18.91 63.99 19.11 505.18 ;
      RECT 18.91 505.38 19.11 510.01 ;
      RECT 18.31 35.31 18.91 35.51 ;
      RECT 18.66 28.03 18.86 28.77 ;
      RECT 18.51 30.13 18.83 30.73 ;
      RECT 18.51 42.75 18.83 43.35 ;
      RECT 18.51 65.96 18.71 510.01 ;
      RECT 17.01 6.24 18.41 6.84 ;
      RECT 18.11 505.38 18.31 510.01 ;
      RECT 17.57 12.98 18.17 13.18 ;
      RECT 17.71 505.38 17.91 510.01 ;
      RECT 17.11 35.31 17.71 35.51 ;
      RECT 17.19 30.13 17.51 30.73 ;
      RECT 17.19 42.75 17.51 43.35 ;
      RECT 9.11 28.15 17.31 28.75 ;
      RECT 16.51 59.37 17.15 59.97 ;
      RECT 16.91 63.99 17.11 505.18 ;
      RECT 16.91 505.38 17.11 510.01 ;
      RECT 16.51 505.38 16.71 510.01 ;
      RECT 14.61 6.24 16.59 6.84 ;
      RECT 15.91 35.31 16.51 35.51 ;
      RECT 16.11 30.13 16.43 30.73 ;
      RECT 16.11 42.75 16.43 43.35 ;
      RECT 15.71 505.38 15.91 510.01 ;
      RECT 15.31 505.38 15.51 510.01 ;
      RECT 14.71 35.31 15.31 35.51 ;
      RECT 14.79 30.13 15.11 30.73 ;
      RECT 14.79 42.75 15.11 43.35 ;
      RECT 14.91 65.96 15.11 510.01 ;
      RECT 14.07 59.37 14.71 59.97 ;
      RECT 14.51 505.38 14.71 510.01 ;
      RECT 14.11 63.99 14.31 505.18 ;
      RECT 14.11 505.38 14.31 510.01 ;
      RECT 12.21 6.24 14.19 6.84 ;
      RECT 13.51 35.31 14.11 35.51 ;
      RECT 13.71 30.13 14.03 30.73 ;
      RECT 13.71 42.75 14.03 43.35 ;
      RECT 12.51 15.51 13.91 15.71 ;
      RECT 13.71 65.96 13.91 510.01 ;
      RECT 13.31 505.38 13.51 510.01 ;
      RECT 12.91 505.38 13.11 510.01 ;
      RECT 12.31 35.31 12.91 35.51 ;
      RECT 12.39 30.13 12.71 30.73 ;
      RECT 12.39 42.75 12.71 43.35 ;
      RECT 11.71 59.37 12.35 59.97 ;
      RECT 12.11 63.99 12.31 505.18 ;
      RECT 12.11 505.38 12.31 510.01 ;
      RECT 11.71 505.38 11.91 510.01 ;
      RECT 9.81 6.24 11.79 6.84 ;
      RECT 11.11 35.31 11.71 35.51 ;
      RECT 11.31 30.13 11.63 30.73 ;
      RECT 11.31 42.75 11.63 43.35 ;
      RECT 10.91 505.38 11.11 510.01 ;
      RECT 10.51 505.38 10.71 510.01 ;
      RECT 9.91 35.31 10.51 35.51 ;
      RECT 9.99 30.13 10.31 30.73 ;
      RECT 9.99 42.75 10.31 43.35 ;
      RECT 10.11 65.96 10.31 510.01 ;
      RECT 9.27 59.37 9.91 59.97 ;
      RECT 9.71 505.38 9.91 510.01 ;
      RECT 9.31 63.99 9.51 505.18 ;
      RECT 9.31 505.38 9.51 510.01 ;
      RECT 7.41 6.24 9.41 6.84 ;
      RECT 8.71 35.31 9.31 35.51 ;
      RECT 8.91 30.13 9.23 30.73 ;
      RECT 8.91 42.75 9.23 43.35 ;
      RECT 8.91 65.96 9.11 510.01 ;
      RECT 8.51 505.38 8.71 510.01 ;
      RECT 7.71 68.76 7.91 70.2 ;
      RECT 7.71 70.4 7.91 71.16 ;
      RECT 7.71 71.36 7.91 72.12 ;
      RECT 7.71 72.32 7.91 73.6 ;
      RECT 7.71 73.8 7.91 74.56 ;
      RECT 7.71 74.76 7.91 75.52 ;
      RECT 7.71 75.72 7.91 77 ;
      RECT 7.71 77.2 7.91 77.96 ;
      RECT 7.71 78.16 7.91 78.92 ;
      RECT 7.71 79.12 7.91 80.4 ;
      RECT 7.71 80.6 7.91 81.36 ;
      RECT 7.71 81.56 7.91 82.32 ;
      RECT 7.71 82.52 7.91 83.8 ;
      RECT 7.71 84 7.91 84.76 ;
      RECT 7.71 84.96 7.91 85.72 ;
      RECT 7.71 85.92 7.91 87.2 ;
      RECT 7.71 87.4 7.91 88.16 ;
      RECT 7.71 88.36 7.91 89.12 ;
      RECT 7.71 89.32 7.91 90.6 ;
      RECT 7.71 90.8 7.91 91.56 ;
      RECT 7.71 91.76 7.91 92.52 ;
      RECT 7.71 92.72 7.91 94 ;
      RECT 7.71 94.2 7.91 94.96 ;
      RECT 7.71 95.16 7.91 95.92 ;
      RECT 7.71 96.12 7.91 97.4 ;
      RECT 7.71 97.6 7.91 98.36 ;
      RECT 7.71 98.56 7.91 99.32 ;
      RECT 7.71 99.52 7.91 100.8 ;
      RECT 7.71 101 7.91 101.76 ;
      RECT 7.71 101.96 7.91 102.72 ;
      RECT 7.71 102.92 7.91 104.2 ;
      RECT 7.71 104.4 7.91 105.16 ;
      RECT 7.71 105.36 7.91 106.12 ;
      RECT 7.71 106.32 7.91 107.6 ;
      RECT 7.71 107.8 7.91 108.56 ;
      RECT 7.71 108.76 7.91 109.52 ;
      RECT 7.71 109.72 7.91 111 ;
      RECT 7.71 111.2 7.91 111.96 ;
      RECT 7.71 112.16 7.91 112.92 ;
      RECT 7.71 113.12 7.91 114.4 ;
      RECT 7.71 114.6 7.91 115.36 ;
      RECT 7.71 115.56 7.91 116.32 ;
      RECT 7.71 116.52 7.91 117.8 ;
      RECT 7.71 118 7.91 118.76 ;
      RECT 7.71 118.96 7.91 119.72 ;
      RECT 7.71 119.92 7.91 121.2 ;
      RECT 7.71 121.4 7.91 122.16 ;
      RECT 7.71 122.36 7.91 123.12 ;
      RECT 7.71 123.32 7.91 124.6 ;
      RECT 7.71 124.8 7.91 125.56 ;
      RECT 7.71 125.76 7.91 126.52 ;
      RECT 7.71 126.72 7.91 128 ;
      RECT 7.71 128.2 7.91 128.96 ;
      RECT 7.71 129.16 7.91 129.92 ;
      RECT 7.71 130.12 7.91 131.4 ;
      RECT 7.71 131.6 7.91 132.36 ;
      RECT 7.71 132.56 7.91 133.32 ;
      RECT 7.71 133.52 7.91 134.8 ;
      RECT 7.71 135 7.91 135.76 ;
      RECT 7.71 135.96 7.91 136.72 ;
      RECT 7.71 136.92 7.91 138.2 ;
      RECT 7.71 138.4 7.91 139.16 ;
      RECT 7.71 139.36 7.91 140.12 ;
      RECT 7.71 140.32 7.91 141.6 ;
      RECT 7.71 141.8 7.91 142.56 ;
      RECT 7.71 142.76 7.91 143.52 ;
      RECT 7.71 143.72 7.91 145 ;
      RECT 7.71 145.2 7.91 145.96 ;
      RECT 7.71 146.16 7.91 146.92 ;
      RECT 7.71 147.12 7.91 148.4 ;
      RECT 7.71 148.6 7.91 149.36 ;
      RECT 7.71 149.56 7.91 150.32 ;
      RECT 7.71 150.52 7.91 151.8 ;
      RECT 7.71 152 7.91 152.76 ;
      RECT 7.71 152.96 7.91 153.72 ;
      RECT 7.71 153.92 7.91 155.2 ;
      RECT 7.71 155.4 7.91 156.16 ;
      RECT 7.71 156.36 7.91 157.12 ;
      RECT 7.71 157.32 7.91 158.6 ;
      RECT 7.71 158.8 7.91 159.56 ;
      RECT 7.71 159.76 7.91 160.52 ;
      RECT 7.71 160.72 7.91 162 ;
      RECT 7.71 162.2 7.91 162.96 ;
      RECT 7.71 163.16 7.91 163.92 ;
      RECT 7.71 164.12 7.91 165.4 ;
      RECT 7.71 165.6 7.91 166.36 ;
      RECT 7.71 166.56 7.91 167.32 ;
      RECT 7.71 167.52 7.91 168.8 ;
      RECT 7.71 169 7.91 169.76 ;
      RECT 7.71 169.96 7.91 170.72 ;
      RECT 7.71 170.92 7.91 172.2 ;
      RECT 7.71 172.4 7.91 173.16 ;
      RECT 7.71 173.36 7.91 174.12 ;
      RECT 7.71 174.32 7.91 175.6 ;
      RECT 7.71 175.8 7.91 176.56 ;
      RECT 7.71 176.76 7.91 177.52 ;
      RECT 7.71 177.72 7.91 179 ;
      RECT 7.71 179.2 7.91 179.96 ;
      RECT 7.71 180.16 7.91 180.92 ;
      RECT 7.71 181.12 7.91 182.4 ;
      RECT 7.71 182.6 7.91 183.36 ;
      RECT 7.71 183.56 7.91 184.32 ;
      RECT 7.71 184.52 7.91 185.8 ;
      RECT 7.71 186 7.91 186.76 ;
      RECT 7.71 186.96 7.91 187.72 ;
      RECT 7.71 187.92 7.91 189.2 ;
      RECT 7.71 189.4 7.91 190.16 ;
      RECT 7.71 190.36 7.91 191.12 ;
      RECT 7.71 191.32 7.91 192.6 ;
      RECT 7.71 192.8 7.91 193.56 ;
      RECT 7.71 193.76 7.91 194.52 ;
      RECT 7.71 194.72 7.91 196 ;
      RECT 7.71 196.2 7.91 196.96 ;
      RECT 7.71 197.16 7.91 197.92 ;
      RECT 7.71 198.12 7.91 199.4 ;
      RECT 7.71 199.6 7.91 200.36 ;
      RECT 7.71 200.56 7.91 201.32 ;
      RECT 7.71 201.52 7.91 202.8 ;
      RECT 7.71 203 7.91 203.76 ;
      RECT 7.71 203.96 7.91 204.72 ;
      RECT 7.71 204.92 7.91 206.2 ;
      RECT 7.71 206.4 7.91 207.16 ;
      RECT 7.71 207.36 7.91 208.12 ;
      RECT 7.71 208.32 7.91 209.6 ;
      RECT 7.71 209.8 7.91 210.56 ;
      RECT 7.71 210.76 7.91 211.52 ;
      RECT 7.71 211.72 7.91 213 ;
      RECT 7.71 213.2 7.91 213.96 ;
      RECT 7.71 214.16 7.91 214.92 ;
      RECT 7.71 215.12 7.91 216.4 ;
      RECT 7.71 216.6 7.91 217.36 ;
      RECT 7.71 217.56 7.91 218.32 ;
      RECT 7.71 218.52 7.91 219.8 ;
      RECT 7.71 220 7.91 220.76 ;
      RECT 7.71 220.96 7.91 221.72 ;
      RECT 7.71 221.92 7.91 223.2 ;
      RECT 7.71 223.4 7.91 224.16 ;
      RECT 7.71 224.36 7.91 225.12 ;
      RECT 7.71 225.32 7.91 226.6 ;
      RECT 7.71 226.8 7.91 227.56 ;
      RECT 7.71 227.76 7.91 228.52 ;
      RECT 7.71 228.72 7.91 230 ;
      RECT 7.71 230.2 7.91 230.96 ;
      RECT 7.71 231.16 7.91 231.92 ;
      RECT 7.71 232.12 7.91 233.4 ;
      RECT 7.71 233.6 7.91 234.36 ;
      RECT 7.71 234.56 7.91 235.32 ;
      RECT 7.71 235.52 7.91 236.8 ;
      RECT 7.71 237 7.91 237.76 ;
      RECT 7.71 237.96 7.91 238.72 ;
      RECT 7.71 238.92 7.91 240.2 ;
      RECT 7.71 240.4 7.91 241.16 ;
      RECT 7.71 241.36 7.91 242.12 ;
      RECT 7.71 242.32 7.91 243.6 ;
      RECT 7.71 243.8 7.91 244.56 ;
      RECT 7.71 244.76 7.91 245.52 ;
      RECT 7.71 245.72 7.91 247 ;
      RECT 7.71 247.2 7.91 247.96 ;
      RECT 7.71 248.16 7.91 248.92 ;
      RECT 7.71 249.12 7.91 250.4 ;
      RECT 7.71 250.6 7.91 251.36 ;
      RECT 7.71 251.56 7.91 252.32 ;
      RECT 7.71 252.52 7.91 253.8 ;
      RECT 7.71 254 7.91 254.76 ;
      RECT 7.71 254.96 7.91 255.72 ;
      RECT 7.71 255.92 7.91 257.2 ;
      RECT 7.71 257.4 7.91 258.16 ;
      RECT 7.71 258.36 7.91 259.12 ;
      RECT 7.71 259.32 7.91 260.6 ;
      RECT 7.71 260.8 7.91 261.56 ;
      RECT 7.71 261.76 7.91 262.52 ;
      RECT 7.71 262.72 7.91 264 ;
      RECT 7.71 264.2 7.91 264.96 ;
      RECT 7.71 265.16 7.91 265.92 ;
      RECT 7.71 266.12 7.91 267.4 ;
      RECT 7.71 267.6 7.91 268.36 ;
      RECT 7.71 268.56 7.91 269.32 ;
      RECT 7.71 269.52 7.91 270.8 ;
      RECT 7.71 271 7.91 271.76 ;
      RECT 7.71 271.96 7.91 272.72 ;
      RECT 7.71 272.92 7.91 274.2 ;
      RECT 7.71 274.4 7.91 275.16 ;
      RECT 7.71 275.36 7.91 276.12 ;
      RECT 7.71 276.32 7.91 277.6 ;
      RECT 7.71 277.8 7.91 278.56 ;
      RECT 7.71 278.76 7.91 279.52 ;
      RECT 7.71 279.72 7.91 281 ;
      RECT 7.71 281.2 7.91 281.96 ;
      RECT 7.71 282.16 7.91 282.92 ;
      RECT 7.71 283.12 7.91 284.4 ;
      RECT 7.71 284.6 7.91 285.36 ;
      RECT 7.71 285.56 7.91 286.32 ;
      RECT 7.71 286.52 7.91 287.8 ;
      RECT 7.71 288 7.91 288.76 ;
      RECT 7.71 288.96 7.91 289.72 ;
      RECT 7.71 289.92 7.91 291.2 ;
      RECT 7.71 291.4 7.91 292.16 ;
      RECT 7.71 292.36 7.91 293.12 ;
      RECT 7.71 293.32 7.91 294.6 ;
      RECT 7.71 294.8 7.91 295.56 ;
      RECT 7.71 295.76 7.91 296.52 ;
      RECT 7.71 296.72 7.91 298 ;
      RECT 7.71 298.2 7.91 298.96 ;
      RECT 7.71 299.16 7.91 299.92 ;
      RECT 7.71 300.12 7.91 301.4 ;
      RECT 7.71 301.6 7.91 302.36 ;
      RECT 7.71 302.56 7.91 303.32 ;
      RECT 7.71 303.52 7.91 304.8 ;
      RECT 7.71 305 7.91 305.76 ;
      RECT 7.71 305.96 7.91 306.72 ;
      RECT 7.71 306.92 7.91 308.2 ;
      RECT 7.71 308.4 7.91 309.16 ;
      RECT 7.71 309.36 7.91 310.12 ;
      RECT 7.71 310.32 7.91 311.6 ;
      RECT 7.71 311.8 7.91 312.56 ;
      RECT 7.71 312.76 7.91 313.52 ;
      RECT 7.71 313.72 7.91 315 ;
      RECT 7.71 315.2 7.91 315.96 ;
      RECT 7.71 316.16 7.91 316.92 ;
      RECT 7.71 317.12 7.91 318.4 ;
      RECT 7.71 318.6 7.91 319.36 ;
      RECT 7.71 319.56 7.91 320.32 ;
      RECT 7.71 320.52 7.91 321.8 ;
      RECT 7.71 322 7.91 322.76 ;
      RECT 7.71 322.96 7.91 323.72 ;
      RECT 7.71 323.92 7.91 325.2 ;
      RECT 7.71 325.4 7.91 326.16 ;
      RECT 7.71 326.36 7.91 327.12 ;
      RECT 7.71 327.32 7.91 328.6 ;
      RECT 7.71 328.8 7.91 329.56 ;
      RECT 7.71 329.76 7.91 330.52 ;
      RECT 7.71 330.72 7.91 332 ;
      RECT 7.71 332.2 7.91 332.96 ;
      RECT 7.71 333.16 7.91 333.92 ;
      RECT 7.71 334.12 7.91 335.4 ;
      RECT 7.71 335.6 7.91 336.36 ;
      RECT 7.71 336.56 7.91 337.32 ;
      RECT 7.71 337.52 7.91 338.8 ;
      RECT 7.71 339 7.91 339.76 ;
      RECT 7.71 339.96 7.91 340.72 ;
      RECT 7.71 340.92 7.91 342.2 ;
      RECT 7.71 342.4 7.91 343.16 ;
      RECT 7.71 343.36 7.91 344.12 ;
      RECT 7.71 344.32 7.91 345.6 ;
      RECT 7.71 345.8 7.91 346.56 ;
      RECT 7.71 346.76 7.91 347.52 ;
      RECT 7.71 347.72 7.91 349 ;
      RECT 7.71 349.2 7.91 349.96 ;
      RECT 7.71 350.16 7.91 350.92 ;
      RECT 7.71 351.12 7.91 352.4 ;
      RECT 7.71 352.6 7.91 353.36 ;
      RECT 7.71 353.56 7.91 354.32 ;
      RECT 7.71 354.52 7.91 355.8 ;
      RECT 7.71 356 7.91 356.76 ;
      RECT 7.71 356.96 7.91 357.72 ;
      RECT 7.71 357.92 7.91 359.2 ;
      RECT 7.71 359.4 7.91 360.16 ;
      RECT 7.71 360.36 7.91 361.12 ;
      RECT 7.71 361.32 7.91 362.6 ;
      RECT 7.71 362.8 7.91 363.56 ;
      RECT 7.71 363.76 7.91 364.52 ;
      RECT 7.71 364.72 7.91 366 ;
      RECT 7.71 366.2 7.91 366.96 ;
      RECT 7.71 367.16 7.91 367.92 ;
      RECT 7.71 368.12 7.91 369.4 ;
      RECT 7.71 369.6 7.91 370.36 ;
      RECT 7.71 370.56 7.91 371.32 ;
      RECT 7.71 371.52 7.91 372.8 ;
      RECT 7.71 373 7.91 373.76 ;
      RECT 7.71 373.96 7.91 374.72 ;
      RECT 7.71 374.92 7.91 376.2 ;
      RECT 7.71 376.4 7.91 377.16 ;
      RECT 7.71 377.36 7.91 378.12 ;
      RECT 7.71 378.32 7.91 379.6 ;
      RECT 7.71 379.8 7.91 380.56 ;
      RECT 7.71 380.76 7.91 381.52 ;
      RECT 7.71 381.72 7.91 383 ;
      RECT 7.71 383.2 7.91 383.96 ;
      RECT 7.71 384.16 7.91 384.92 ;
      RECT 7.71 385.12 7.91 386.4 ;
      RECT 7.71 386.6 7.91 387.36 ;
      RECT 7.71 387.56 7.91 388.32 ;
      RECT 7.71 388.52 7.91 389.8 ;
      RECT 7.71 390 7.91 390.76 ;
      RECT 7.71 390.96 7.91 391.72 ;
      RECT 7.71 391.92 7.91 393.2 ;
      RECT 7.71 393.4 7.91 394.16 ;
      RECT 7.71 394.36 7.91 395.12 ;
      RECT 7.71 395.32 7.91 396.6 ;
      RECT 7.71 396.8 7.91 397.56 ;
      RECT 7.71 397.76 7.91 398.52 ;
      RECT 7.71 398.72 7.91 400 ;
      RECT 7.71 400.2 7.91 400.96 ;
      RECT 7.71 401.16 7.91 401.92 ;
      RECT 7.71 402.12 7.91 403.4 ;
      RECT 7.71 403.6 7.91 404.36 ;
      RECT 7.71 404.56 7.91 405.32 ;
      RECT 7.71 405.52 7.91 406.8 ;
      RECT 7.71 407 7.91 407.76 ;
      RECT 7.71 407.96 7.91 408.72 ;
      RECT 7.71 408.92 7.91 410.2 ;
      RECT 7.71 410.4 7.91 411.16 ;
      RECT 7.71 411.36 7.91 412.12 ;
      RECT 7.71 412.32 7.91 413.6 ;
      RECT 7.71 413.8 7.91 414.56 ;
      RECT 7.71 414.76 7.91 415.52 ;
      RECT 7.71 415.72 7.91 417 ;
      RECT 7.71 417.2 7.91 417.96 ;
      RECT 7.71 418.16 7.91 418.92 ;
      RECT 7.71 419.12 7.91 420.4 ;
      RECT 7.71 420.6 7.91 421.36 ;
      RECT 7.71 421.56 7.91 422.32 ;
      RECT 7.71 422.52 7.91 423.8 ;
      RECT 7.71 424 7.91 424.76 ;
      RECT 7.71 424.96 7.91 425.72 ;
      RECT 7.71 425.92 7.91 427.2 ;
      RECT 7.71 427.4 7.91 428.16 ;
      RECT 7.71 428.36 7.91 429.12 ;
      RECT 7.71 429.32 7.91 430.6 ;
      RECT 7.71 430.8 7.91 431.56 ;
      RECT 7.71 431.76 7.91 432.52 ;
      RECT 7.71 432.72 7.91 434 ;
      RECT 7.71 434.2 7.91 434.96 ;
      RECT 7.71 435.16 7.91 435.92 ;
      RECT 7.71 436.12 7.91 437.4 ;
      RECT 7.71 437.6 7.91 438.36 ;
      RECT 7.71 438.56 7.91 439.32 ;
      RECT 7.71 439.52 7.91 440.8 ;
      RECT 7.71 441 7.91 441.76 ;
      RECT 7.71 441.96 7.91 442.72 ;
      RECT 7.71 442.92 7.91 444.2 ;
      RECT 7.71 444.4 7.91 445.16 ;
      RECT 7.71 445.36 7.91 446.12 ;
      RECT 7.71 446.32 7.91 447.6 ;
      RECT 7.71 447.8 7.91 448.56 ;
      RECT 7.71 448.76 7.91 449.52 ;
      RECT 7.71 449.72 7.91 451 ;
      RECT 7.71 451.2 7.91 451.96 ;
      RECT 7.71 452.16 7.91 452.92 ;
      RECT 7.71 453.12 7.91 454.4 ;
      RECT 7.71 454.6 7.91 455.36 ;
      RECT 7.71 455.56 7.91 456.32 ;
      RECT 7.71 456.52 7.91 457.8 ;
      RECT 7.71 458 7.91 458.76 ;
      RECT 7.71 458.96 7.91 459.72 ;
      RECT 7.71 459.92 7.91 461.2 ;
      RECT 7.71 461.4 7.91 462.16 ;
      RECT 7.71 462.36 7.91 463.12 ;
      RECT 7.71 463.32 7.91 464.6 ;
      RECT 7.71 464.8 7.91 465.56 ;
      RECT 7.71 465.76 7.91 466.52 ;
      RECT 7.71 466.72 7.91 468 ;
      RECT 7.71 468.2 7.91 468.96 ;
      RECT 7.71 469.16 7.91 469.92 ;
      RECT 7.71 470.12 7.91 471.4 ;
      RECT 7.71 471.6 7.91 472.36 ;
      RECT 7.71 472.56 7.91 473.32 ;
      RECT 7.71 473.52 7.91 474.8 ;
      RECT 7.71 475 7.91 475.76 ;
      RECT 7.71 475.96 7.91 476.72 ;
      RECT 7.71 476.92 7.91 478.2 ;
      RECT 7.71 478.4 7.91 479.16 ;
      RECT 7.71 479.36 7.91 480.12 ;
      RECT 7.71 480.32 7.91 481.6 ;
      RECT 7.71 481.8 7.91 482.56 ;
      RECT 7.71 482.76 7.91 483.52 ;
      RECT 7.71 483.72 7.91 485 ;
      RECT 7.71 485.2 7.91 485.96 ;
      RECT 7.71 486.16 7.91 486.92 ;
      RECT 7.71 487.12 7.91 488.4 ;
      RECT 7.71 488.6 7.91 489.36 ;
      RECT 7.71 489.56 7.91 490.32 ;
      RECT 7.71 490.52 7.91 491.8 ;
      RECT 7.71 492 7.91 492.76 ;
      RECT 7.71 492.96 7.91 493.72 ;
      RECT 7.71 493.92 7.91 495.2 ;
      RECT 7.71 495.4 7.91 496.16 ;
      RECT 7.71 496.36 7.91 497.12 ;
      RECT 7.71 497.32 7.91 498.6 ;
      RECT 7.71 498.8 7.91 499.56 ;
      RECT 7.71 499.76 7.91 500.52 ;
      RECT 7.71 500.72 7.91 502 ;
      RECT 7.71 502.2 7.91 502.96 ;
      RECT 7.71 503.16 7.91 503.92 ;
      RECT 7.71 504.12 7.91 506.44 ;
      RECT 7.71 506.64 7.91 507.4 ;
      RECT 7.71 507.6 7.91 508.36 ;
      RECT 7.71 508.56 7.91 510 ;
      RECT 6.24 12.64 6.84 13.74 ;
      RECT 6.24 69.16 6.84 69.96 ;
      RECT 6.24 72.56 6.84 73.36 ;
      RECT 6.24 75.96 6.84 76.76 ;
      RECT 6.24 79.36 6.84 80.16 ;
      RECT 6.24 82.76 6.84 83.56 ;
      RECT 6.24 86.16 6.84 86.96 ;
      RECT 6.24 89.56 6.84 90.36 ;
      RECT 6.24 92.96 6.84 93.76 ;
      RECT 6.24 96.36 6.84 97.16 ;
      RECT 6.24 99.76 6.84 100.56 ;
      RECT 6.24 103.16 6.84 103.96 ;
      RECT 6.24 106.56 6.84 107.36 ;
      RECT 6.24 109.96 6.84 110.76 ;
      RECT 6.24 113.36 6.84 114.16 ;
      RECT 6.24 116.76 6.84 117.56 ;
      RECT 6.24 120.16 6.84 120.96 ;
      RECT 6.24 123.56 6.84 124.36 ;
      RECT 6.24 126.96 6.84 127.76 ;
      RECT 6.24 130.36 6.84 131.16 ;
      RECT 6.24 133.76 6.84 134.56 ;
      RECT 6.24 137.16 6.84 137.96 ;
      RECT 6.24 140.56 6.84 141.36 ;
      RECT 6.24 143.96 6.84 144.76 ;
      RECT 6.24 147.36 6.84 148.16 ;
      RECT 6.24 150.76 6.84 151.56 ;
      RECT 6.24 154.16 6.84 154.96 ;
      RECT 6.24 157.56 6.84 158.36 ;
      RECT 6.24 160.96 6.84 161.76 ;
      RECT 6.24 164.36 6.84 165.16 ;
      RECT 6.24 167.76 6.84 168.56 ;
      RECT 6.24 171.16 6.84 171.96 ;
      RECT 6.24 174.56 6.84 175.36 ;
      RECT 6.24 177.96 6.84 178.76 ;
      RECT 6.24 181.36 6.84 182.16 ;
      RECT 6.24 184.76 6.84 185.56 ;
      RECT 6.24 188.16 6.84 188.96 ;
      RECT 6.24 191.56 6.84 192.36 ;
      RECT 6.24 194.96 6.84 195.76 ;
      RECT 6.24 198.36 6.84 199.16 ;
      RECT 6.24 201.76 6.84 202.56 ;
      RECT 6.24 205.16 6.84 205.96 ;
      RECT 6.24 208.56 6.84 209.36 ;
      RECT 6.24 211.96 6.84 212.76 ;
      RECT 6.24 215.36 6.84 216.16 ;
      RECT 6.24 218.76 6.84 219.56 ;
      RECT 6.24 222.16 6.84 222.96 ;
      RECT 6.24 225.56 6.84 226.36 ;
      RECT 6.24 228.96 6.84 229.76 ;
      RECT 6.24 232.36 6.84 233.16 ;
      RECT 6.24 235.76 6.84 236.56 ;
      RECT 6.24 239.16 6.84 239.96 ;
      RECT 6.24 242.56 6.84 243.36 ;
      RECT 6.24 245.96 6.84 246.76 ;
      RECT 6.24 249.36 6.84 250.16 ;
      RECT 6.24 252.76 6.84 253.56 ;
      RECT 6.24 256.16 6.84 256.96 ;
      RECT 6.24 259.56 6.84 260.36 ;
      RECT 6.24 262.96 6.84 263.76 ;
      RECT 6.24 266.36 6.84 267.16 ;
      RECT 6.24 269.76 6.84 270.56 ;
      RECT 6.24 273.16 6.84 273.96 ;
      RECT 6.24 276.56 6.84 277.36 ;
      RECT 6.24 279.96 6.84 280.76 ;
      RECT 6.24 283.36 6.84 284.16 ;
      RECT 6.24 286.76 6.84 287.56 ;
      RECT 6.24 290.16 6.84 290.96 ;
      RECT 6.24 293.56 6.84 294.36 ;
      RECT 6.24 296.96 6.84 297.76 ;
      RECT 6.24 300.36 6.84 301.16 ;
      RECT 6.24 303.76 6.84 304.56 ;
      RECT 6.24 307.16 6.84 307.96 ;
      RECT 6.24 310.56 6.84 311.36 ;
      RECT 6.24 313.96 6.84 314.76 ;
      RECT 6.24 317.36 6.84 318.16 ;
      RECT 6.24 320.76 6.84 321.56 ;
      RECT 6.24 324.16 6.84 324.96 ;
      RECT 6.24 327.56 6.84 328.36 ;
      RECT 6.24 330.96 6.84 331.76 ;
      RECT 6.24 334.36 6.84 335.16 ;
      RECT 6.24 337.76 6.84 338.56 ;
      RECT 6.24 341.16 6.84 341.96 ;
      RECT 6.24 344.56 6.84 345.36 ;
      RECT 6.24 347.96 6.84 348.76 ;
      RECT 6.24 351.36 6.84 352.16 ;
      RECT 6.24 354.76 6.84 355.56 ;
      RECT 6.24 358.16 6.84 358.96 ;
      RECT 6.24 361.56 6.84 362.36 ;
      RECT 6.24 364.96 6.84 365.76 ;
      RECT 6.24 368.36 6.84 369.16 ;
      RECT 6.24 371.76 6.84 372.56 ;
      RECT 6.24 375.16 6.84 375.96 ;
      RECT 6.24 378.56 6.84 379.36 ;
      RECT 6.24 381.96 6.84 382.76 ;
      RECT 6.24 385.36 6.84 386.16 ;
      RECT 6.24 388.76 6.84 389.56 ;
      RECT 6.24 392.16 6.84 392.96 ;
      RECT 6.24 395.56 6.84 396.36 ;
      RECT 6.24 398.96 6.84 399.76 ;
      RECT 6.24 402.36 6.84 403.16 ;
      RECT 6.24 405.76 6.84 406.56 ;
      RECT 6.24 409.16 6.84 409.96 ;
      RECT 6.24 412.56 6.84 413.36 ;
      RECT 6.24 415.96 6.84 416.76 ;
      RECT 6.24 419.36 6.84 420.16 ;
      RECT 6.24 422.76 6.84 423.56 ;
      RECT 6.24 426.16 6.84 426.96 ;
      RECT 6.24 429.56 6.84 430.36 ;
      RECT 6.24 432.96 6.84 433.76 ;
      RECT 6.24 436.36 6.84 437.16 ;
      RECT 6.24 439.76 6.84 440.56 ;
      RECT 6.24 443.16 6.84 443.96 ;
      RECT 6.24 446.56 6.84 447.36 ;
      RECT 6.24 449.96 6.84 450.76 ;
      RECT 6.24 453.36 6.84 454.16 ;
      RECT 6.24 456.76 6.84 457.56 ;
      RECT 6.24 460.16 6.84 460.96 ;
      RECT 6.24 463.56 6.84 464.36 ;
      RECT 6.24 466.96 6.84 467.76 ;
      RECT 6.24 470.36 6.84 471.16 ;
      RECT 6.24 473.76 6.84 474.56 ;
      RECT 6.24 477.16 6.84 477.96 ;
      RECT 6.24 480.56 6.84 481.36 ;
      RECT 6.24 483.96 6.84 484.76 ;
      RECT 6.24 487.36 6.84 488.16 ;
      RECT 6.24 490.76 6.84 491.56 ;
      RECT 6.24 494.16 6.84 494.96 ;
      RECT 6.24 497.56 6.84 498.36 ;
      RECT 6.24 500.96 6.84 501.76 ;
      RECT 6.24 504.36 6.84 505.16 ;
      RECT 6.24 505.6 6.84 506 ;
      RECT 6.24 509 6.84 509.8 ;
    LAYER M3 ;
      RECT 228.79 509 230.79 510.94 ;
      RECT 223.99 509 225.99 510.94 ;
      RECT 219.19 509 221.19 510.94 ;
      RECT 214.39 509 216.39 510.94 ;
      RECT 209.59 509 211.59 510.94 ;
      RECT 204.79 509 206.79 510.94 ;
      RECT 199.99 509 201.99 510.94 ;
      RECT 195.19 509 197.19 510.94 ;
      RECT 189.19 509 191.19 510.94 ;
      RECT 184.39 509 186.39 510.94 ;
      RECT 179.59 509 181.59 510.94 ;
      RECT 174.79 509 176.79 510.94 ;
      RECT 169.99 509 171.99 510.94 ;
      RECT 165.19 509 167.19 510.94 ;
      RECT 160.39 509 162.39 510.94 ;
      RECT 155.59 509 157.59 510.94 ;
      RECT 148.01 32.39 149.33 510.94 ;
      RECT 233.76 509 240.6 509.8 ;
      RECT 148.01 509.2 152.7 509.6 ;
      RECT 152.3 509 240.6 509.4 ;
      RECT 148.01 505.6 240.6 506 ;
      RECT 233.76 504.36 240.6 505.16 ;
      RECT 148.01 504.56 240.6 504.96 ;
      RECT 233.76 500.96 240.6 501.76 ;
      RECT 148.01 501.16 240.6 501.56 ;
      RECT 233.76 497.56 240.6 498.36 ;
      RECT 148.01 497.76 240.6 498.16 ;
      RECT 233.76 494.16 240.6 494.96 ;
      RECT 148.01 494.36 240.6 494.76 ;
      RECT 233.76 490.76 240.6 491.56 ;
      RECT 148.01 490.96 240.6 491.36 ;
      RECT 233.76 487.36 240.6 488.16 ;
      RECT 148.01 487.56 240.6 487.96 ;
      RECT 233.76 483.96 240.6 484.76 ;
      RECT 148.01 484.16 240.6 484.56 ;
      RECT 233.76 480.56 240.6 481.36 ;
      RECT 148.01 480.76 240.6 481.16 ;
      RECT 233.76 477.16 240.6 477.96 ;
      RECT 148.01 477.36 240.6 477.76 ;
      RECT 233.76 473.76 240.6 474.56 ;
      RECT 148.01 473.96 240.6 474.36 ;
      RECT 233.76 470.36 240.6 471.16 ;
      RECT 148.01 470.56 240.6 470.96 ;
      RECT 233.76 466.96 240.6 467.76 ;
      RECT 148.01 467.16 240.6 467.56 ;
      RECT 233.76 463.56 240.6 464.36 ;
      RECT 148.01 463.76 240.6 464.16 ;
      RECT 233.76 460.16 240.6 460.96 ;
      RECT 148.01 460.36 240.6 460.76 ;
      RECT 233.76 456.76 240.6 457.56 ;
      RECT 148.01 456.96 240.6 457.36 ;
      RECT 233.76 453.36 240.6 454.16 ;
      RECT 148.01 453.56 240.6 453.96 ;
      RECT 233.76 449.96 240.6 450.76 ;
      RECT 148.01 450.16 240.6 450.56 ;
      RECT 233.76 446.56 240.6 447.36 ;
      RECT 148.01 446.76 240.6 447.16 ;
      RECT 233.76 443.16 240.6 443.96 ;
      RECT 148.01 443.36 240.6 443.76 ;
      RECT 233.76 439.76 240.6 440.56 ;
      RECT 148.01 439.96 240.6 440.36 ;
      RECT 233.76 436.36 240.6 437.16 ;
      RECT 148.01 436.56 240.6 436.96 ;
      RECT 233.76 432.96 240.6 433.76 ;
      RECT 148.01 433.16 240.6 433.56 ;
      RECT 233.76 429.56 240.6 430.36 ;
      RECT 148.01 429.76 240.6 430.16 ;
      RECT 233.76 426.16 240.6 426.96 ;
      RECT 148.01 426.36 240.6 426.76 ;
      RECT 233.76 422.76 240.6 423.56 ;
      RECT 148.01 422.96 240.6 423.36 ;
      RECT 233.76 419.36 240.6 420.16 ;
      RECT 148.01 419.56 240.6 419.96 ;
      RECT 233.76 415.96 240.6 416.76 ;
      RECT 148.01 416.16 240.6 416.56 ;
      RECT 233.76 412.56 240.6 413.36 ;
      RECT 148.01 412.76 240.6 413.16 ;
      RECT 233.76 409.16 240.6 409.96 ;
      RECT 148.01 409.36 240.6 409.76 ;
      RECT 233.76 405.76 240.6 406.56 ;
      RECT 148.01 405.96 240.6 406.36 ;
      RECT 233.76 402.36 240.6 403.16 ;
      RECT 148.01 402.56 240.6 402.96 ;
      RECT 233.76 398.96 240.6 399.76 ;
      RECT 148.01 399.16 240.6 399.56 ;
      RECT 233.76 395.56 240.6 396.36 ;
      RECT 148.01 395.76 240.6 396.16 ;
      RECT 233.76 392.16 240.6 392.96 ;
      RECT 148.01 392.36 240.6 392.76 ;
      RECT 233.76 388.76 240.6 389.56 ;
      RECT 148.01 388.96 240.6 389.36 ;
      RECT 233.76 385.36 240.6 386.16 ;
      RECT 148.01 385.56 240.6 385.96 ;
      RECT 233.76 381.96 240.6 382.76 ;
      RECT 148.01 382.16 240.6 382.56 ;
      RECT 233.76 378.56 240.6 379.36 ;
      RECT 148.01 378.76 240.6 379.16 ;
      RECT 233.76 375.16 240.6 375.96 ;
      RECT 148.01 375.36 240.6 375.76 ;
      RECT 233.76 371.76 240.6 372.56 ;
      RECT 148.01 371.96 240.6 372.36 ;
      RECT 233.76 368.36 240.6 369.16 ;
      RECT 148.01 368.56 240.6 368.96 ;
      RECT 233.76 364.96 240.6 365.76 ;
      RECT 148.01 365.16 240.6 365.56 ;
      RECT 233.76 361.56 240.6 362.36 ;
      RECT 148.01 361.76 240.6 362.16 ;
      RECT 233.76 358.16 240.6 358.96 ;
      RECT 148.01 358.36 240.6 358.76 ;
      RECT 233.76 354.76 240.6 355.56 ;
      RECT 148.01 354.96 240.6 355.36 ;
      RECT 233.76 351.36 240.6 352.16 ;
      RECT 148.01 351.56 240.6 351.96 ;
      RECT 233.76 347.96 240.6 348.76 ;
      RECT 148.01 348.16 240.6 348.56 ;
      RECT 233.76 344.56 240.6 345.36 ;
      RECT 148.01 344.76 240.6 345.16 ;
      RECT 233.76 341.16 240.6 341.96 ;
      RECT 148.01 341.36 240.6 341.76 ;
      RECT 233.76 337.76 240.6 338.56 ;
      RECT 148.01 337.96 240.6 338.36 ;
      RECT 233.76 334.36 240.6 335.16 ;
      RECT 148.01 334.56 240.6 334.96 ;
      RECT 233.76 330.96 240.6 331.76 ;
      RECT 148.01 331.16 240.6 331.56 ;
      RECT 233.76 327.56 240.6 328.36 ;
      RECT 148.01 327.76 240.6 328.16 ;
      RECT 233.76 324.16 240.6 324.96 ;
      RECT 148.01 324.36 240.6 324.76 ;
      RECT 233.76 320.76 240.6 321.56 ;
      RECT 148.01 320.96 240.6 321.36 ;
      RECT 233.76 317.36 240.6 318.16 ;
      RECT 148.01 317.56 240.6 317.96 ;
      RECT 233.76 313.96 240.6 314.76 ;
      RECT 148.01 314.16 240.6 314.56 ;
      RECT 233.76 310.56 240.6 311.36 ;
      RECT 148.01 310.76 240.6 311.16 ;
      RECT 233.76 307.16 240.6 307.96 ;
      RECT 148.01 307.36 240.6 307.76 ;
      RECT 233.76 303.76 240.6 304.56 ;
      RECT 148.01 303.96 240.6 304.36 ;
      RECT 233.76 300.36 240.6 301.16 ;
      RECT 148.01 300.56 240.6 300.96 ;
      RECT 233.76 296.96 240.6 297.76 ;
      RECT 148.01 297.16 240.6 297.56 ;
      RECT 233.76 293.56 240.6 294.36 ;
      RECT 148.01 293.76 240.6 294.16 ;
      RECT 233.76 290.16 240.6 290.96 ;
      RECT 148.01 290.36 240.6 290.76 ;
      RECT 233.76 286.76 240.6 287.56 ;
      RECT 148.01 286.96 240.6 287.36 ;
      RECT 233.76 283.36 240.6 284.16 ;
      RECT 148.01 283.56 240.6 283.96 ;
      RECT 233.76 279.96 240.6 280.76 ;
      RECT 148.01 280.16 240.6 280.56 ;
      RECT 233.76 276.56 240.6 277.36 ;
      RECT 148.01 276.76 240.6 277.16 ;
      RECT 233.76 273.16 240.6 273.96 ;
      RECT 148.01 273.36 240.6 273.76 ;
      RECT 233.76 269.76 240.6 270.56 ;
      RECT 148.01 269.96 240.6 270.36 ;
      RECT 233.76 266.36 240.6 267.16 ;
      RECT 148.01 266.56 240.6 266.96 ;
      RECT 233.76 262.96 240.6 263.76 ;
      RECT 148.01 263.16 240.6 263.56 ;
      RECT 233.76 259.56 240.6 260.36 ;
      RECT 148.01 259.76 240.6 260.16 ;
      RECT 233.76 256.16 240.6 256.96 ;
      RECT 148.01 256.36 240.6 256.76 ;
      RECT 233.76 252.76 240.6 253.56 ;
      RECT 148.01 252.96 240.6 253.36 ;
      RECT 233.76 249.36 240.6 250.16 ;
      RECT 148.01 249.56 240.6 249.96 ;
      RECT 233.76 245.96 240.6 246.76 ;
      RECT 148.01 246.16 240.6 246.56 ;
      RECT 233.76 242.56 240.6 243.36 ;
      RECT 148.01 242.76 240.6 243.16 ;
      RECT 233.76 239.16 240.6 239.96 ;
      RECT 148.01 239.36 240.6 239.76 ;
      RECT 233.76 235.76 240.6 236.56 ;
      RECT 148.01 235.96 240.6 236.36 ;
      RECT 233.76 232.36 240.6 233.16 ;
      RECT 148.01 232.56 240.6 232.96 ;
      RECT 233.76 228.96 240.6 229.76 ;
      RECT 148.01 229.16 240.6 229.56 ;
      RECT 233.76 225.56 240.6 226.36 ;
      RECT 148.01 225.76 240.6 226.16 ;
      RECT 233.76 222.16 240.6 222.96 ;
      RECT 148.01 222.36 240.6 222.76 ;
      RECT 233.76 218.76 240.6 219.56 ;
      RECT 148.01 218.96 240.6 219.36 ;
      RECT 233.76 215.36 240.6 216.16 ;
      RECT 148.01 215.56 240.6 215.96 ;
      RECT 233.76 211.96 240.6 212.76 ;
      RECT 148.01 212.16 240.6 212.56 ;
      RECT 233.76 208.56 240.6 209.36 ;
      RECT 148.01 208.76 240.6 209.16 ;
      RECT 233.76 205.16 240.6 205.96 ;
      RECT 148.01 205.36 240.6 205.76 ;
      RECT 233.76 201.76 240.6 202.56 ;
      RECT 148.01 201.96 240.6 202.36 ;
      RECT 233.76 198.36 240.6 199.16 ;
      RECT 148.01 198.56 240.6 198.96 ;
      RECT 233.76 194.96 240.6 195.76 ;
      RECT 148.01 195.16 240.6 195.56 ;
      RECT 233.76 191.56 240.6 192.36 ;
      RECT 148.01 191.76 240.6 192.16 ;
      RECT 233.76 188.16 240.6 188.96 ;
      RECT 148.01 188.36 240.6 188.76 ;
      RECT 233.76 184.76 240.6 185.56 ;
      RECT 148.01 184.96 240.6 185.36 ;
      RECT 233.76 181.36 240.6 182.16 ;
      RECT 148.01 181.56 240.6 181.96 ;
      RECT 233.76 177.96 240.6 178.76 ;
      RECT 148.01 178.16 240.6 178.56 ;
      RECT 233.76 174.56 240.6 175.36 ;
      RECT 148.01 174.76 240.6 175.16 ;
      RECT 233.76 171.16 240.6 171.96 ;
      RECT 148.01 171.36 240.6 171.76 ;
      RECT 233.76 167.76 240.6 168.56 ;
      RECT 148.01 167.96 240.6 168.36 ;
      RECT 233.76 164.36 240.6 165.16 ;
      RECT 148.01 164.56 240.6 164.96 ;
      RECT 233.76 160.96 240.6 161.76 ;
      RECT 148.01 161.16 240.6 161.56 ;
      RECT 233.76 157.56 240.6 158.36 ;
      RECT 148.01 157.76 240.6 158.16 ;
      RECT 233.76 154.16 240.6 154.96 ;
      RECT 148.01 154.36 240.6 154.76 ;
      RECT 233.76 150.76 240.6 151.56 ;
      RECT 148.01 150.96 240.6 151.36 ;
      RECT 233.76 147.36 240.6 148.16 ;
      RECT 148.01 147.56 240.6 147.96 ;
      RECT 233.76 143.96 240.6 144.76 ;
      RECT 148.01 144.16 240.6 144.56 ;
      RECT 233.76 140.56 240.6 141.36 ;
      RECT 148.01 140.76 240.6 141.16 ;
      RECT 233.76 137.16 240.6 137.96 ;
      RECT 148.01 137.36 240.6 137.76 ;
      RECT 233.76 133.76 240.6 134.56 ;
      RECT 148.01 133.96 240.6 134.36 ;
      RECT 233.76 130.36 240.6 131.16 ;
      RECT 148.01 130.56 240.6 130.96 ;
      RECT 233.76 126.96 240.6 127.76 ;
      RECT 148.01 127.16 240.6 127.56 ;
      RECT 233.76 123.56 240.6 124.36 ;
      RECT 148.01 123.76 240.6 124.16 ;
      RECT 233.76 120.16 240.6 120.96 ;
      RECT 148.01 120.36 240.6 120.76 ;
      RECT 233.76 116.76 240.6 117.56 ;
      RECT 148.01 116.96 240.6 117.36 ;
      RECT 233.76 113.36 240.6 114.16 ;
      RECT 148.01 113.56 240.6 113.96 ;
      RECT 233.76 109.96 240.6 110.76 ;
      RECT 148.01 110.16 240.6 110.56 ;
      RECT 233.76 106.56 240.6 107.36 ;
      RECT 148.01 106.76 240.6 107.16 ;
      RECT 233.76 103.16 240.6 103.96 ;
      RECT 148.01 103.36 240.6 103.76 ;
      RECT 233.76 99.76 240.6 100.56 ;
      RECT 148.01 99.96 240.6 100.36 ;
      RECT 233.76 96.36 240.6 97.16 ;
      RECT 148.01 96.56 240.6 96.96 ;
      RECT 233.76 92.96 240.6 93.76 ;
      RECT 148.01 93.16 240.6 93.56 ;
      RECT 233.76 89.56 240.6 90.36 ;
      RECT 148.01 89.76 240.6 90.16 ;
      RECT 233.76 86.16 240.6 86.96 ;
      RECT 148.01 86.36 240.6 86.76 ;
      RECT 233.76 82.76 240.6 83.56 ;
      RECT 148.01 82.96 240.6 83.36 ;
      RECT 233.76 79.36 240.6 80.16 ;
      RECT 148.01 79.56 240.6 79.96 ;
      RECT 233.76 75.96 240.6 76.76 ;
      RECT 148.01 76.16 240.6 76.56 ;
      RECT 233.76 72.56 240.6 73.36 ;
      RECT 148.01 72.76 240.6 73.16 ;
      RECT 233.76 69.16 240.6 69.96 ;
      RECT 148.01 69.36 240.6 69.76 ;
      RECT 148.47 6.24 148.87 510.94 ;
      RECT 148.01 6.24 148.87 8.59 ;
      RECT 230.29 67.59 233.39 68.59 ;
      RECT 232.79 6.24 233.19 68.59 ;
      RECT 231.99 6.24 232.39 68.59 ;
      RECT 232.79 54.22 237.48 55.22 ;
      RECT 232.79 41.29 237.48 42.29 ;
      RECT 232.79 39.44 237.48 40.44 ;
      RECT 230.69 37.61 231.29 37.81 ;
      RECT 230.69 28.55 230.89 37.81 ;
      RECT 231.09 28.55 231.29 37.41 ;
      RECT 232.79 32.98 237.48 33.98 ;
      RECT 232.79 31.13 237.48 32.13 ;
      RECT 230.69 28.55 232.39 28.75 ;
      RECT 231.29 28.15 232.39 28.75 ;
      RECT 232.79 21.41 237.48 22.21 ;
      RECT 232.79 12.64 237.48 13.74 ;
      RECT 231.19 6.24 233.19 6.84 ;
      RECT 233.76 70.86 237.48 71.66 ;
      RECT 149.73 71.06 237.48 71.46 ;
      RECT 233.76 74.26 237.48 75.06 ;
      RECT 149.73 74.46 237.48 74.86 ;
      RECT 233.76 77.66 237.48 78.46 ;
      RECT 149.73 77.86 237.48 78.26 ;
      RECT 233.76 81.06 237.48 81.86 ;
      RECT 149.73 81.26 237.48 81.66 ;
      RECT 233.76 84.46 237.48 85.26 ;
      RECT 149.73 84.66 237.48 85.06 ;
      RECT 233.76 87.86 237.48 88.66 ;
      RECT 149.73 88.06 237.48 88.46 ;
      RECT 233.76 91.26 237.48 92.06 ;
      RECT 149.73 91.46 237.48 91.86 ;
      RECT 233.76 94.66 237.48 95.46 ;
      RECT 149.73 94.86 237.48 95.26 ;
      RECT 233.76 98.06 237.48 98.86 ;
      RECT 149.73 98.26 237.48 98.66 ;
      RECT 233.76 101.46 237.48 102.26 ;
      RECT 149.73 101.66 237.48 102.06 ;
      RECT 233.76 104.86 237.48 105.66 ;
      RECT 149.73 105.06 237.48 105.46 ;
      RECT 233.76 108.26 237.48 109.06 ;
      RECT 149.73 108.46 237.48 108.86 ;
      RECT 233.76 111.66 237.48 112.46 ;
      RECT 149.73 111.86 237.48 112.26 ;
      RECT 233.76 115.06 237.48 115.86 ;
      RECT 149.73 115.26 237.48 115.66 ;
      RECT 233.76 118.46 237.48 119.26 ;
      RECT 149.73 118.66 237.48 119.06 ;
      RECT 233.76 121.86 237.48 122.66 ;
      RECT 149.73 122.06 237.48 122.46 ;
      RECT 233.76 125.26 237.48 126.06 ;
      RECT 149.73 125.46 237.48 125.86 ;
      RECT 233.76 128.66 237.48 129.46 ;
      RECT 149.73 128.86 237.48 129.26 ;
      RECT 233.76 132.06 237.48 132.86 ;
      RECT 149.73 132.26 237.48 132.66 ;
      RECT 233.76 135.46 237.48 136.26 ;
      RECT 149.73 135.66 237.48 136.06 ;
      RECT 233.76 138.86 237.48 139.66 ;
      RECT 149.73 139.06 237.48 139.46 ;
      RECT 233.76 142.26 237.48 143.06 ;
      RECT 149.73 142.46 237.48 142.86 ;
      RECT 233.76 145.66 237.48 146.46 ;
      RECT 149.73 145.86 237.48 146.26 ;
      RECT 233.76 149.06 237.48 149.86 ;
      RECT 149.73 149.26 237.48 149.66 ;
      RECT 233.76 152.46 237.48 153.26 ;
      RECT 149.73 152.66 237.48 153.06 ;
      RECT 233.76 155.86 237.48 156.66 ;
      RECT 149.73 156.06 237.48 156.46 ;
      RECT 233.76 159.26 237.48 160.06 ;
      RECT 149.73 159.46 237.48 159.86 ;
      RECT 233.76 162.66 237.48 163.46 ;
      RECT 149.73 162.86 237.48 163.26 ;
      RECT 233.76 166.06 237.48 166.86 ;
      RECT 149.73 166.26 237.48 166.66 ;
      RECT 233.76 169.46 237.48 170.26 ;
      RECT 149.73 169.66 237.48 170.06 ;
      RECT 233.76 172.86 237.48 173.66 ;
      RECT 149.73 173.06 237.48 173.46 ;
      RECT 233.76 176.26 237.48 177.06 ;
      RECT 149.73 176.46 237.48 176.86 ;
      RECT 233.76 179.66 237.48 180.46 ;
      RECT 149.73 179.86 237.48 180.26 ;
      RECT 233.76 183.06 237.48 183.86 ;
      RECT 149.73 183.26 237.48 183.66 ;
      RECT 233.76 186.46 237.48 187.26 ;
      RECT 149.73 186.66 237.48 187.06 ;
      RECT 233.76 189.86 237.48 190.66 ;
      RECT 149.73 190.06 237.48 190.46 ;
      RECT 233.76 193.26 237.48 194.06 ;
      RECT 149.73 193.46 237.48 193.86 ;
      RECT 233.76 196.66 237.48 197.46 ;
      RECT 149.73 196.86 237.48 197.26 ;
      RECT 233.76 200.06 237.48 200.86 ;
      RECT 149.73 200.26 237.48 200.66 ;
      RECT 233.76 203.46 237.48 204.26 ;
      RECT 149.73 203.66 237.48 204.06 ;
      RECT 233.76 206.86 237.48 207.66 ;
      RECT 149.73 207.06 237.48 207.46 ;
      RECT 233.76 210.26 237.48 211.06 ;
      RECT 149.73 210.46 237.48 210.86 ;
      RECT 233.76 213.66 237.48 214.46 ;
      RECT 149.73 213.86 237.48 214.26 ;
      RECT 233.76 217.06 237.48 217.86 ;
      RECT 149.73 217.26 237.48 217.66 ;
      RECT 233.76 220.46 237.48 221.26 ;
      RECT 149.73 220.66 237.48 221.06 ;
      RECT 233.76 223.86 237.48 224.66 ;
      RECT 149.73 224.06 237.48 224.46 ;
      RECT 233.76 227.26 237.48 228.06 ;
      RECT 149.73 227.46 237.48 227.86 ;
      RECT 233.76 230.66 237.48 231.46 ;
      RECT 149.73 230.86 237.48 231.26 ;
      RECT 233.76 234.06 237.48 234.86 ;
      RECT 149.73 234.26 237.48 234.66 ;
      RECT 233.76 237.46 237.48 238.26 ;
      RECT 149.73 237.66 237.48 238.06 ;
      RECT 233.76 240.86 237.48 241.66 ;
      RECT 149.73 241.06 237.48 241.46 ;
      RECT 233.76 244.26 237.48 245.06 ;
      RECT 149.73 244.46 237.48 244.86 ;
      RECT 233.76 247.66 237.48 248.46 ;
      RECT 149.73 247.86 237.48 248.26 ;
      RECT 233.76 251.06 237.48 251.86 ;
      RECT 149.73 251.26 237.48 251.66 ;
      RECT 233.76 254.46 237.48 255.26 ;
      RECT 149.73 254.66 237.48 255.06 ;
      RECT 233.76 257.86 237.48 258.66 ;
      RECT 149.73 258.06 237.48 258.46 ;
      RECT 233.76 261.26 237.48 262.06 ;
      RECT 149.73 261.46 237.48 261.86 ;
      RECT 233.76 264.66 237.48 265.46 ;
      RECT 149.73 264.86 237.48 265.26 ;
      RECT 233.76 268.06 237.48 268.86 ;
      RECT 149.73 268.26 237.48 268.66 ;
      RECT 233.76 271.46 237.48 272.26 ;
      RECT 149.73 271.66 237.48 272.06 ;
      RECT 233.76 274.86 237.48 275.66 ;
      RECT 149.73 275.06 237.48 275.46 ;
      RECT 233.76 278.26 237.48 279.06 ;
      RECT 149.73 278.46 237.48 278.86 ;
      RECT 233.76 281.66 237.48 282.46 ;
      RECT 149.73 281.86 237.48 282.26 ;
      RECT 233.76 285.06 237.48 285.86 ;
      RECT 149.73 285.26 237.48 285.66 ;
      RECT 233.76 288.46 237.48 289.26 ;
      RECT 149.73 288.66 237.48 289.06 ;
      RECT 233.76 291.86 237.48 292.66 ;
      RECT 149.73 292.06 237.48 292.46 ;
      RECT 233.76 295.26 237.48 296.06 ;
      RECT 149.73 295.46 237.48 295.86 ;
      RECT 233.76 298.66 237.48 299.46 ;
      RECT 149.73 298.86 237.48 299.26 ;
      RECT 233.76 302.06 237.48 302.86 ;
      RECT 149.73 302.26 237.48 302.66 ;
      RECT 233.76 305.46 237.48 306.26 ;
      RECT 149.73 305.66 237.48 306.06 ;
      RECT 233.76 308.86 237.48 309.66 ;
      RECT 149.73 309.06 237.48 309.46 ;
      RECT 233.76 312.26 237.48 313.06 ;
      RECT 149.73 312.46 237.48 312.86 ;
      RECT 233.76 315.66 237.48 316.46 ;
      RECT 149.73 315.86 237.48 316.26 ;
      RECT 233.76 319.06 237.48 319.86 ;
      RECT 149.73 319.26 237.48 319.66 ;
      RECT 233.76 322.46 237.48 323.26 ;
      RECT 149.73 322.66 237.48 323.06 ;
      RECT 233.76 325.86 237.48 326.66 ;
      RECT 149.73 326.06 237.48 326.46 ;
      RECT 233.76 329.26 237.48 330.06 ;
      RECT 149.73 329.46 237.48 329.86 ;
      RECT 233.76 332.66 237.48 333.46 ;
      RECT 149.73 332.86 237.48 333.26 ;
      RECT 233.76 336.06 237.48 336.86 ;
      RECT 149.73 336.26 237.48 336.66 ;
      RECT 233.76 339.46 237.48 340.26 ;
      RECT 149.73 339.66 237.48 340.06 ;
      RECT 233.76 342.86 237.48 343.66 ;
      RECT 149.73 343.06 237.48 343.46 ;
      RECT 233.76 346.26 237.48 347.06 ;
      RECT 149.73 346.46 237.48 346.86 ;
      RECT 233.76 349.66 237.48 350.46 ;
      RECT 149.73 349.86 237.48 350.26 ;
      RECT 233.76 353.06 237.48 353.86 ;
      RECT 149.73 353.26 237.48 353.66 ;
      RECT 233.76 356.46 237.48 357.26 ;
      RECT 149.73 356.66 237.48 357.06 ;
      RECT 233.76 359.86 237.48 360.66 ;
      RECT 149.73 360.06 237.48 360.46 ;
      RECT 233.76 363.26 237.48 364.06 ;
      RECT 149.73 363.46 237.48 363.86 ;
      RECT 233.76 366.66 237.48 367.46 ;
      RECT 149.73 366.86 237.48 367.26 ;
      RECT 233.76 370.06 237.48 370.86 ;
      RECT 149.73 370.26 237.48 370.66 ;
      RECT 233.76 373.46 237.48 374.26 ;
      RECT 149.73 373.66 237.48 374.06 ;
      RECT 233.76 376.86 237.48 377.66 ;
      RECT 149.73 377.06 237.48 377.46 ;
      RECT 233.76 380.26 237.48 381.06 ;
      RECT 149.73 380.46 237.48 380.86 ;
      RECT 233.76 383.66 237.48 384.46 ;
      RECT 149.73 383.86 237.48 384.26 ;
      RECT 233.76 387.06 237.48 387.86 ;
      RECT 149.73 387.26 237.48 387.66 ;
      RECT 233.76 390.46 237.48 391.26 ;
      RECT 149.73 390.66 237.48 391.06 ;
      RECT 233.76 393.86 237.48 394.66 ;
      RECT 149.73 394.06 237.48 394.46 ;
      RECT 233.76 397.26 237.48 398.06 ;
      RECT 149.73 397.46 237.48 397.86 ;
      RECT 233.76 400.66 237.48 401.46 ;
      RECT 149.73 400.86 237.48 401.26 ;
      RECT 233.76 404.06 237.48 404.86 ;
      RECT 149.73 404.26 237.48 404.66 ;
      RECT 233.76 407.46 237.48 408.26 ;
      RECT 149.73 407.66 237.48 408.06 ;
      RECT 233.76 410.86 237.48 411.66 ;
      RECT 149.73 411.06 237.48 411.46 ;
      RECT 233.76 414.26 237.48 415.06 ;
      RECT 149.73 414.46 237.48 414.86 ;
      RECT 233.76 417.66 237.48 418.46 ;
      RECT 149.73 417.86 237.48 418.26 ;
      RECT 233.76 421.06 237.48 421.86 ;
      RECT 149.73 421.26 237.48 421.66 ;
      RECT 233.76 424.46 237.48 425.26 ;
      RECT 149.73 424.66 237.48 425.06 ;
      RECT 233.76 427.86 237.48 428.66 ;
      RECT 149.73 428.06 237.48 428.46 ;
      RECT 233.76 431.26 237.48 432.06 ;
      RECT 149.73 431.46 237.48 431.86 ;
      RECT 233.76 434.66 237.48 435.46 ;
      RECT 149.73 434.86 237.48 435.26 ;
      RECT 233.76 438.06 237.48 438.86 ;
      RECT 149.73 438.26 237.48 438.66 ;
      RECT 233.76 441.46 237.48 442.26 ;
      RECT 149.73 441.66 237.48 442.06 ;
      RECT 233.76 444.86 237.48 445.66 ;
      RECT 149.73 445.06 237.48 445.46 ;
      RECT 233.76 448.26 237.48 449.06 ;
      RECT 149.73 448.46 237.48 448.86 ;
      RECT 233.76 451.66 237.48 452.46 ;
      RECT 149.73 451.86 237.48 452.26 ;
      RECT 233.76 455.06 237.48 455.86 ;
      RECT 149.73 455.26 237.48 455.66 ;
      RECT 233.76 458.46 237.48 459.26 ;
      RECT 149.73 458.66 237.48 459.06 ;
      RECT 233.76 461.86 237.48 462.66 ;
      RECT 149.73 462.06 237.48 462.46 ;
      RECT 233.76 465.26 237.48 466.06 ;
      RECT 149.73 465.46 237.48 465.86 ;
      RECT 233.76 468.66 237.48 469.46 ;
      RECT 149.73 468.86 237.48 469.26 ;
      RECT 233.76 472.06 237.48 472.86 ;
      RECT 149.73 472.26 237.48 472.66 ;
      RECT 233.76 475.46 237.48 476.26 ;
      RECT 149.73 475.66 237.48 476.06 ;
      RECT 233.76 478.86 237.48 479.66 ;
      RECT 149.73 479.06 237.48 479.46 ;
      RECT 233.76 482.26 237.48 483.06 ;
      RECT 149.73 482.46 237.48 482.86 ;
      RECT 233.76 485.66 237.48 486.46 ;
      RECT 149.73 485.86 237.48 486.26 ;
      RECT 233.76 489.06 237.48 489.86 ;
      RECT 149.73 489.26 237.48 489.66 ;
      RECT 233.76 492.46 237.48 493.26 ;
      RECT 149.73 492.66 237.48 493.06 ;
      RECT 233.76 495.86 237.48 496.66 ;
      RECT 149.73 496.06 237.48 496.46 ;
      RECT 233.76 499.26 237.48 500.06 ;
      RECT 149.73 499.46 237.48 499.86 ;
      RECT 233.76 502.66 237.48 503.46 ;
      RECT 149.73 502.86 237.48 503.26 ;
      RECT 195.41 508.1 237.48 508.6 ;
      RECT 232.89 506.6 237.48 508.6 ;
      RECT 195.41 506.4 195.91 508.6 ;
      RECT 195.41 507.3 237.48 507.7 ;
      RECT 195.41 506.4 233.4 506.9 ;
      RECT 232.39 510.34 233.19 510.94 ;
      RECT 231.19 510.34 231.99 510.94 ;
      RECT 231.19 510.34 233.39 510.74 ;
      RECT 231.09 38.01 231.29 65.45 ;
      RECT 231.09 38.01 231.69 38.21 ;
      RECT 231.49 30.13 231.69 38.21 ;
      RECT 229.59 27.82 229.99 68.59 ;
      RECT 227.89 65.96 231.69 66.96 ;
      RECT 229.99 6.24 230.73 28.22 ;
      RECT 228.81 6.24 230.73 18.31 ;
      RECT 228.81 6.24 230.79 7.44 ;
      RECT 230.69 38.01 230.89 65.05 ;
      RECT 230.29 38.01 230.89 38.21 ;
      RECT 230.29 30.13 230.49 38.21 ;
      RECT 228.69 38.01 228.89 65.05 ;
      RECT 228.69 38.01 229.29 38.21 ;
      RECT 229.09 30.13 229.29 38.21 ;
      RECT 225.49 67.59 229.29 68.59 ;
      RECT 227.19 28.15 227.59 68.59 ;
      RECT 228.29 37.61 228.89 37.81 ;
      RECT 228.69 28.75 228.89 37.81 ;
      RECT 228.29 28.15 228.49 37.41 ;
      RECT 228.29 28.75 228.89 28.95 ;
      RECT 228.29 38.01 228.49 65.45 ;
      RECT 227.89 38.01 228.49 38.21 ;
      RECT 227.89 30.13 228.09 38.21 ;
      RECT 226.69 6.24 228.09 25.07 ;
      RECT 226.41 6.24 228.39 7.44 ;
      RECT 227.59 510.34 228.39 510.94 ;
      RECT 226.39 510.34 227.19 510.94 ;
      RECT 226.39 510.34 228.39 510.74 ;
      RECT 226.29 38.01 226.49 65.45 ;
      RECT 226.29 38.01 226.89 38.21 ;
      RECT 226.69 30.13 226.89 38.21 ;
      RECT 224.79 27.82 225.19 68.59 ;
      RECT 223.09 65.96 226.89 66.96 ;
      RECT 224.05 6.24 224.79 28.22 ;
      RECT 224.05 6.24 225.99 18.31 ;
      RECT 224.01 6.24 225.99 7.44 ;
      RECT 225.89 37.61 226.49 37.81 ;
      RECT 225.89 28.75 226.09 37.81 ;
      RECT 226.29 28.15 226.49 37.41 ;
      RECT 225.89 28.75 226.49 28.95 ;
      RECT 225.89 38.01 226.09 65.05 ;
      RECT 225.49 38.01 226.09 38.21 ;
      RECT 225.49 30.13 225.69 38.21 ;
      RECT 223.89 38.01 224.09 65.05 ;
      RECT 223.89 38.01 224.49 38.21 ;
      RECT 224.29 30.13 224.49 38.21 ;
      RECT 220.69 67.59 224.49 68.59 ;
      RECT 222.39 6.24 222.79 68.59 ;
      RECT 223.49 37.61 224.09 37.81 ;
      RECT 223.89 28.55 224.09 37.81 ;
      RECT 221.09 37.61 221.69 37.81 ;
      RECT 221.09 28.55 221.29 37.81 ;
      RECT 223.49 28.55 223.69 37.41 ;
      RECT 221.49 28.55 221.69 37.41 ;
      RECT 221.49 28.55 222.79 28.95 ;
      RECT 221.09 28.55 224.09 28.75 ;
      RECT 222.39 28.15 223.49 28.75 ;
      RECT 221.99 9.34 222.79 9.54 ;
      RECT 221.59 6.24 223.59 6.84 ;
      RECT 223.49 38.01 223.69 65.45 ;
      RECT 223.09 38.01 223.69 38.21 ;
      RECT 223.09 30.13 223.29 38.21 ;
      RECT 222.79 510.34 223.59 510.94 ;
      RECT 221.59 510.34 222.39 510.94 ;
      RECT 221.59 510.34 223.59 510.74 ;
      RECT 221.49 38.01 221.69 65.45 ;
      RECT 221.49 38.01 222.09 38.21 ;
      RECT 221.89 30.13 222.09 38.21 ;
      RECT 219.99 27.82 220.39 68.59 ;
      RECT 218.29 65.96 222.09 66.96 ;
      RECT 219.99 27.82 221.13 28.22 ;
      RECT 220.93 7.54 221.13 28.22 ;
      RECT 220.39 7.54 221.13 20.81 ;
      RECT 219.99 6.24 220.79 8.24 ;
      RECT 219.21 6.24 221.19 6.84 ;
      RECT 221.74 25.29 221.94 28.35 ;
      RECT 221.53 25.29 221.94 25.49 ;
      RECT 221.53 21.25 221.73 25.49 ;
      RECT 221.09 38.01 221.29 65.05 ;
      RECT 220.69 38.01 221.29 38.21 ;
      RECT 220.69 30.13 220.89 38.21 ;
      RECT 219.59 27.42 219.79 28.57 ;
      RECT 219.59 27.42 220.73 27.62 ;
      RECT 220.53 21.01 220.73 27.62 ;
      RECT 219.99 21.01 220.73 21.21 ;
      RECT 219.99 18.71 220.19 21.21 ;
      RECT 218.69 37.61 219.29 37.81 ;
      RECT 219.09 27.02 219.29 37.81 ;
      RECT 219.09 27.02 220.33 27.22 ;
      RECT 220.13 21.41 220.33 27.22 ;
      RECT 219.59 21.41 220.33 21.61 ;
      RECT 219.59 12.98 219.79 21.61 ;
      RECT 219.73 21.81 219.93 23.85 ;
      RECT 219.19 21.81 219.93 22.01 ;
      RECT 219.19 20.73 219.39 22.01 ;
      RECT 219.09 38.01 219.29 65.05 ;
      RECT 219.09 38.01 219.69 38.21 ;
      RECT 219.49 30.13 219.69 38.21 ;
      RECT 215.89 67.59 219.69 68.59 ;
      RECT 217.59 26.07 217.99 68.59 ;
      RECT 217.09 26.07 217.99 28.61 ;
      RECT 217.09 26.07 218.49 28.6 ;
      RECT 216.43 26.07 219.15 26.27 ;
      RECT 218.95 24.87 219.15 26.27 ;
      RECT 216.43 24.87 216.63 26.27 ;
      RECT 216.43 24.87 219.15 25.07 ;
      RECT 217.09 14.44 218.49 25.07 ;
      RECT 217.59 6.24 217.99 25.07 ;
      RECT 217.29 6.24 218.79 6.84 ;
      RECT 218.69 38.01 218.89 65.45 ;
      RECT 218.29 38.01 218.89 38.21 ;
      RECT 218.29 30.13 218.49 38.21 ;
      RECT 217.99 510.34 218.79 510.94 ;
      RECT 216.79 510.34 217.59 510.94 ;
      RECT 216.79 510.34 218.79 510.74 ;
      RECT 216.29 37.61 216.89 37.81 ;
      RECT 216.29 27.02 216.49 37.81 ;
      RECT 215.25 27.02 216.49 27.22 ;
      RECT 215.25 21.41 215.45 27.22 ;
      RECT 215.25 21.41 215.99 21.61 ;
      RECT 215.79 19.42 215.99 21.61 ;
      RECT 215.79 19.42 216.59 19.62 ;
      RECT 216.39 13.78 216.59 19.62 ;
      RECT 216.39 13.78 217.39 13.98 ;
      RECT 217.19 8.94 217.39 13.98 ;
      RECT 216.69 38.01 216.89 65.45 ;
      RECT 216.69 38.01 217.29 38.21 ;
      RECT 217.09 30.13 217.29 38.21 ;
      RECT 215.19 27.82 215.59 68.59 ;
      RECT 213.49 65.96 217.29 66.96 ;
      RECT 214.45 27.82 215.59 28.22 ;
      RECT 214.45 7.54 214.65 28.22 ;
      RECT 214.45 16.1 215.19 20.81 ;
      RECT 214.05 14.76 214.79 16.84 ;
      RECT 214.45 7.54 215.19 15.5 ;
      RECT 214.89 6.24 215.69 8.24 ;
      RECT 214.89 6.24 215.89 6.84 ;
      RECT 216.79 8.94 216.99 13.58 ;
      RECT 216.52 8.94 216.99 9.14 ;
      RECT 216.29 38.01 216.49 65.05 ;
      RECT 215.89 38.01 216.49 38.21 ;
      RECT 215.89 30.13 216.09 38.21 ;
      RECT 215.65 21.81 215.85 23.85 ;
      RECT 215.65 21.81 216.39 22.01 ;
      RECT 216.19 20.73 216.39 22.01 ;
      RECT 215.79 27.42 215.99 28.57 ;
      RECT 214.85 27.42 215.99 27.62 ;
      RECT 214.85 21.01 215.05 27.62 ;
      RECT 214.85 21.01 215.59 21.21 ;
      RECT 215.39 15.7 215.59 21.21 ;
      RECT 214.99 15.7 215.59 15.9 ;
      RECT 214.29 38.01 214.49 65.05 ;
      RECT 214.29 38.01 214.89 38.21 ;
      RECT 214.69 30.13 214.89 38.21 ;
      RECT 211.09 67.59 214.89 68.59 ;
      RECT 212.79 6.24 213.19 68.59 ;
      RECT 213.89 37.61 214.49 37.81 ;
      RECT 214.29 28.55 214.49 37.81 ;
      RECT 211.49 37.61 212.09 37.81 ;
      RECT 211.49 28.55 211.69 37.81 ;
      RECT 213.89 28.55 214.09 37.41 ;
      RECT 211.89 28.55 212.09 37.41 ;
      RECT 211.89 28.55 214.09 28.95 ;
      RECT 211.49 28.55 214.49 28.75 ;
      RECT 212.59 6.24 213.39 6.84 ;
      RECT 213.39 9.82 213.59 15.58 ;
      RECT 213.39 9.82 214.09 10.02 ;
      RECT 213.89 7.14 214.09 10.02 ;
      RECT 213.89 38.01 214.09 65.45 ;
      RECT 213.49 38.01 214.09 38.21 ;
      RECT 213.49 30.13 213.69 38.21 ;
      RECT 213.64 25.29 213.84 28.35 ;
      RECT 213.64 25.29 214.05 25.49 ;
      RECT 213.85 21.25 214.05 25.49 ;
      RECT 213.19 510.34 213.99 510.94 ;
      RECT 211.99 510.34 212.79 510.94 ;
      RECT 211.99 510.34 213.99 510.74 ;
      RECT 212.39 9.82 212.59 15.58 ;
      RECT 211.89 9.82 212.59 10.02 ;
      RECT 211.89 7.14 212.09 10.02 ;
      RECT 211.89 38.01 212.09 65.45 ;
      RECT 211.89 38.01 212.49 38.21 ;
      RECT 212.29 30.13 212.49 38.21 ;
      RECT 210.39 27.82 210.79 68.59 ;
      RECT 208.69 65.96 212.49 66.96 ;
      RECT 210.39 27.82 211.53 28.22 ;
      RECT 211.33 7.54 211.53 28.22 ;
      RECT 210.79 16.1 211.53 20.81 ;
      RECT 211.19 14.76 211.93 16.84 ;
      RECT 210.79 7.54 211.53 15.5 ;
      RECT 210.29 6.24 211.09 8.24 ;
      RECT 210.09 6.24 211.09 6.84 ;
      RECT 212.14 25.29 212.34 28.35 ;
      RECT 211.93 25.29 212.34 25.49 ;
      RECT 211.93 21.25 212.13 25.49 ;
      RECT 211.49 38.01 211.69 65.05 ;
      RECT 211.09 38.01 211.69 38.21 ;
      RECT 211.09 30.13 211.29 38.21 ;
      RECT 209.99 27.42 210.19 28.57 ;
      RECT 209.99 27.42 211.13 27.62 ;
      RECT 210.93 21.01 211.13 27.62 ;
      RECT 210.39 21.01 211.13 21.21 ;
      RECT 210.39 15.7 210.59 21.21 ;
      RECT 210.39 15.7 210.99 15.9 ;
      RECT 209.09 37.61 209.69 37.81 ;
      RECT 209.49 27.02 209.69 37.81 ;
      RECT 209.49 27.02 210.73 27.22 ;
      RECT 210.53 21.41 210.73 27.22 ;
      RECT 209.99 21.41 210.73 21.61 ;
      RECT 209.99 19.42 210.19 21.61 ;
      RECT 209.39 19.42 210.19 19.62 ;
      RECT 209.39 13.78 209.59 19.62 ;
      RECT 208.59 13.78 209.59 13.98 ;
      RECT 208.59 8.94 208.79 13.98 ;
      RECT 210.13 21.81 210.33 23.85 ;
      RECT 209.59 21.81 210.33 22.01 ;
      RECT 209.59 20.73 209.79 22.01 ;
      RECT 209.49 38.01 209.69 65.05 ;
      RECT 209.49 38.01 210.09 38.21 ;
      RECT 209.89 30.13 210.09 38.21 ;
      RECT 206.29 67.59 210.09 68.59 ;
      RECT 207.99 26.07 208.39 68.59 ;
      RECT 207.99 26.07 208.89 28.61 ;
      RECT 207.49 26.07 208.89 28.6 ;
      RECT 206.83 26.07 209.55 26.27 ;
      RECT 209.35 24.87 209.55 26.27 ;
      RECT 206.83 24.87 207.03 26.27 ;
      RECT 206.83 24.87 209.55 25.07 ;
      RECT 207.49 14.44 208.89 25.07 ;
      RECT 207.99 6.24 208.39 25.07 ;
      RECT 207.19 6.24 208.69 6.84 ;
      RECT 208.99 8.94 209.19 13.58 ;
      RECT 208.99 8.94 209.46 9.14 ;
      RECT 209.09 38.01 209.29 65.45 ;
      RECT 208.69 38.01 209.29 38.21 ;
      RECT 208.69 30.13 208.89 38.21 ;
      RECT 208.39 510.34 209.19 510.94 ;
      RECT 207.19 510.34 207.99 510.94 ;
      RECT 207.19 510.34 209.19 510.74 ;
      RECT 207.09 38.01 207.29 65.45 ;
      RECT 207.09 38.01 207.69 38.21 ;
      RECT 207.49 30.13 207.69 38.21 ;
      RECT 205.59 27.82 205.99 68.59 ;
      RECT 203.89 65.96 207.69 66.96 ;
      RECT 204.85 27.82 205.99 28.22 ;
      RECT 204.85 7.54 205.05 28.22 ;
      RECT 204.85 7.54 205.59 20.81 ;
      RECT 205.19 6.24 205.99 8.24 ;
      RECT 204.79 6.24 206.76 6.84 ;
      RECT 206.69 37.61 207.29 37.81 ;
      RECT 206.69 27.02 206.89 37.81 ;
      RECT 205.65 27.02 206.89 27.22 ;
      RECT 205.65 21.41 205.85 27.22 ;
      RECT 205.65 21.41 206.39 21.61 ;
      RECT 206.19 12.98 206.39 21.61 ;
      RECT 206.69 38.01 206.89 65.05 ;
      RECT 206.29 38.01 206.89 38.21 ;
      RECT 206.29 30.13 206.49 38.21 ;
      RECT 206.05 21.81 206.25 23.85 ;
      RECT 206.05 21.81 206.79 22.01 ;
      RECT 206.59 20.73 206.79 22.01 ;
      RECT 206.19 27.42 206.39 28.57 ;
      RECT 205.25 27.42 206.39 27.62 ;
      RECT 205.25 21.01 205.45 27.62 ;
      RECT 205.25 21.01 205.99 21.21 ;
      RECT 205.79 18.71 205.99 21.21 ;
      RECT 204.69 38.01 204.89 65.05 ;
      RECT 204.69 38.01 205.29 38.21 ;
      RECT 205.09 30.13 205.29 38.21 ;
      RECT 201.49 67.59 205.29 68.59 ;
      RECT 203.19 6.24 203.59 68.59 ;
      RECT 204.29 37.61 204.89 37.81 ;
      RECT 204.69 28.55 204.89 37.81 ;
      RECT 201.89 37.61 202.49 37.81 ;
      RECT 201.89 28.55 202.09 37.81 ;
      RECT 204.29 28.55 204.49 37.41 ;
      RECT 202.29 28.55 202.49 37.41 ;
      RECT 203.19 28.55 204.49 28.95 ;
      RECT 201.89 28.55 204.89 28.75 ;
      RECT 202.49 28.15 203.59 28.75 ;
      RECT 203.19 9.34 203.99 9.54 ;
      RECT 202.39 6.24 204.39 6.84 ;
      RECT 204.29 38.01 204.49 65.45 ;
      RECT 203.89 38.01 204.49 38.21 ;
      RECT 203.89 30.13 204.09 38.21 ;
      RECT 204.04 25.29 204.24 28.35 ;
      RECT 204.04 25.29 204.45 25.49 ;
      RECT 204.25 21.25 204.45 25.49 ;
      RECT 203.59 510.34 204.39 510.94 ;
      RECT 202.39 510.34 203.19 510.94 ;
      RECT 202.39 510.34 204.39 510.74 ;
      RECT 202.29 38.01 202.49 65.45 ;
      RECT 202.29 38.01 202.89 38.21 ;
      RECT 202.69 30.13 202.89 38.21 ;
      RECT 200.79 27.82 201.19 68.59 ;
      RECT 199.09 65.96 202.89 66.96 ;
      RECT 201.19 6.24 201.93 28.22 ;
      RECT 199.99 6.24 201.93 18.31 ;
      RECT 199.99 6.24 201.97 7.44 ;
      RECT 201.89 38.01 202.09 65.05 ;
      RECT 201.49 38.01 202.09 38.21 ;
      RECT 201.49 30.13 201.69 38.21 ;
      RECT 199.89 38.01 200.09 65.05 ;
      RECT 199.89 38.01 200.49 38.21 ;
      RECT 200.29 30.13 200.49 38.21 ;
      RECT 196.69 67.59 200.49 68.59 ;
      RECT 198.39 28.15 198.79 68.59 ;
      RECT 199.49 37.61 200.09 37.81 ;
      RECT 199.89 28.75 200.09 37.81 ;
      RECT 199.49 28.15 199.69 37.41 ;
      RECT 199.49 28.75 200.09 28.95 ;
      RECT 199.49 38.01 199.69 65.45 ;
      RECT 199.09 38.01 199.69 38.21 ;
      RECT 199.09 30.13 199.29 38.21 ;
      RECT 198.79 510.34 199.59 510.94 ;
      RECT 197.59 510.34 198.39 510.94 ;
      RECT 197.59 510.34 199.59 510.74 ;
      RECT 197.89 6.24 199.29 25.07 ;
      RECT 197.59 6.24 199.57 7.44 ;
      RECT 197.49 38.01 197.69 65.45 ;
      RECT 197.49 38.01 198.09 38.21 ;
      RECT 197.89 30.13 198.09 38.21 ;
      RECT 195.99 27.82 196.39 68.59 ;
      RECT 194.29 65.96 198.09 66.96 ;
      RECT 195.25 6.24 195.99 28.22 ;
      RECT 195.25 6.24 197.17 18.31 ;
      RECT 195.19 6.24 197.17 7.44 ;
      RECT 197.09 37.61 197.69 37.81 ;
      RECT 197.09 28.75 197.29 37.81 ;
      RECT 197.49 28.15 197.69 37.41 ;
      RECT 197.09 28.75 197.69 28.95 ;
      RECT 197.09 38.01 197.29 65.05 ;
      RECT 196.69 38.01 197.29 38.21 ;
      RECT 196.69 30.13 196.89 38.21 ;
      RECT 195.09 38.01 195.29 65.05 ;
      RECT 195.09 38.01 195.69 38.21 ;
      RECT 195.49 30.13 195.69 38.21 ;
      RECT 193.59 67.59 195.69 68.59 ;
      RECT 190.69 67.59 192.79 68.59 ;
      RECT 192.39 6.24 192.79 68.59 ;
      RECT 193.59 6.24 193.99 68.59 ;
      RECT 192.99 7.04 193.39 55.22 ;
      RECT 194.69 37.61 195.29 37.81 ;
      RECT 195.09 28.55 195.29 37.81 ;
      RECT 191.09 37.61 191.69 37.81 ;
      RECT 191.09 28.55 191.29 37.81 ;
      RECT 194.69 28.55 194.89 37.41 ;
      RECT 191.49 28.55 191.69 37.41 ;
      RECT 193.59 28.55 195.29 28.75 ;
      RECT 191.09 28.55 192.79 28.75 ;
      RECT 191.69 28.15 192.79 28.75 ;
      RECT 193.59 28.15 194.69 28.75 ;
      RECT 193.39 6.24 193.99 9.04 ;
      RECT 192.39 6.24 192.99 9.04 ;
      RECT 193.39 6.24 194.79 6.84 ;
      RECT 191.59 6.24 192.99 6.84 ;
      RECT 149.61 508.1 195 508.6 ;
      RECT 194.5 506.4 195 508.6 ;
      RECT 150.13 506.4 195 506.9 ;
      RECT 194.69 38.01 194.89 65.45 ;
      RECT 194.29 38.01 194.89 38.21 ;
      RECT 194.29 30.13 194.49 38.21 ;
      RECT 193.99 510.34 194.79 510.94 ;
      RECT 192.79 510.34 193.59 510.94 ;
      RECT 191.59 510.34 192.39 510.94 ;
      RECT 191.59 510.34 194.79 510.74 ;
      RECT 149.63 507.3 150.03 507.81 ;
      RECT 149.63 507.3 194.09 507.7 ;
      RECT 191.49 38.01 191.69 65.45 ;
      RECT 191.49 38.01 192.09 38.21 ;
      RECT 191.89 30.13 192.09 38.21 ;
      RECT 189.99 27.82 190.39 68.59 ;
      RECT 188.29 65.96 192.09 66.96 ;
      RECT 190.39 6.24 191.13 28.22 ;
      RECT 189.21 6.24 191.13 18.31 ;
      RECT 189.21 6.24 191.19 7.44 ;
      RECT 191.09 38.01 191.29 65.05 ;
      RECT 190.69 38.01 191.29 38.21 ;
      RECT 190.69 30.13 190.89 38.21 ;
      RECT 189.09 38.01 189.29 65.05 ;
      RECT 189.09 38.01 189.69 38.21 ;
      RECT 189.49 30.13 189.69 38.21 ;
      RECT 185.89 67.59 189.69 68.59 ;
      RECT 187.59 28.15 187.99 68.59 ;
      RECT 188.69 37.61 189.29 37.81 ;
      RECT 189.09 28.75 189.29 37.81 ;
      RECT 188.69 28.15 188.89 37.41 ;
      RECT 188.69 28.75 189.29 28.95 ;
      RECT 188.69 38.01 188.89 65.45 ;
      RECT 188.29 38.01 188.89 38.21 ;
      RECT 188.29 30.13 188.49 38.21 ;
      RECT 187.09 6.24 188.49 25.07 ;
      RECT 186.81 6.24 188.79 7.44 ;
      RECT 187.99 510.34 188.79 510.94 ;
      RECT 186.79 510.34 187.59 510.94 ;
      RECT 186.79 510.34 188.79 510.74 ;
      RECT 186.69 38.01 186.89 65.45 ;
      RECT 186.69 38.01 187.29 38.21 ;
      RECT 187.09 30.13 187.29 38.21 ;
      RECT 185.19 27.82 185.59 68.59 ;
      RECT 183.49 65.96 187.29 66.96 ;
      RECT 184.45 6.24 185.19 28.22 ;
      RECT 184.45 6.24 186.39 18.31 ;
      RECT 184.41 6.24 186.39 7.44 ;
      RECT 186.29 37.61 186.89 37.81 ;
      RECT 186.29 28.75 186.49 37.81 ;
      RECT 186.69 28.15 186.89 37.41 ;
      RECT 186.29 28.75 186.89 28.95 ;
      RECT 186.29 38.01 186.49 65.05 ;
      RECT 185.89 38.01 186.49 38.21 ;
      RECT 185.89 30.13 186.09 38.21 ;
      RECT 184.29 38.01 184.49 65.05 ;
      RECT 184.29 38.01 184.89 38.21 ;
      RECT 184.69 30.13 184.89 38.21 ;
      RECT 181.09 67.59 184.89 68.59 ;
      RECT 182.79 6.24 183.19 68.59 ;
      RECT 183.89 37.61 184.49 37.81 ;
      RECT 184.29 28.55 184.49 37.81 ;
      RECT 181.49 37.61 182.09 37.81 ;
      RECT 181.49 28.55 181.69 37.81 ;
      RECT 183.89 28.55 184.09 37.41 ;
      RECT 181.89 28.55 182.09 37.41 ;
      RECT 181.89 28.55 183.19 28.95 ;
      RECT 181.49 28.55 184.49 28.75 ;
      RECT 182.79 28.15 183.89 28.75 ;
      RECT 182.39 9.34 183.19 9.54 ;
      RECT 181.99 6.24 183.99 6.84 ;
      RECT 183.89 38.01 184.09 65.45 ;
      RECT 183.49 38.01 184.09 38.21 ;
      RECT 183.49 30.13 183.69 38.21 ;
      RECT 183.19 510.34 183.99 510.94 ;
      RECT 181.99 510.34 182.79 510.94 ;
      RECT 181.99 510.34 183.99 510.74 ;
      RECT 181.89 38.01 182.09 65.45 ;
      RECT 181.89 38.01 182.49 38.21 ;
      RECT 182.29 30.13 182.49 38.21 ;
      RECT 180.39 27.82 180.79 68.59 ;
      RECT 178.69 65.96 182.49 66.96 ;
      RECT 180.39 27.82 181.53 28.22 ;
      RECT 181.33 7.54 181.53 28.22 ;
      RECT 180.79 7.54 181.53 20.81 ;
      RECT 180.39 6.24 181.19 8.24 ;
      RECT 179.62 6.24 181.59 6.84 ;
      RECT 182.14 25.29 182.34 28.35 ;
      RECT 181.93 25.29 182.34 25.49 ;
      RECT 181.93 21.25 182.13 25.49 ;
      RECT 181.49 38.01 181.69 65.05 ;
      RECT 181.09 38.01 181.69 38.21 ;
      RECT 181.09 30.13 181.29 38.21 ;
      RECT 179.99 27.42 180.19 28.57 ;
      RECT 179.99 27.42 181.13 27.62 ;
      RECT 180.93 21.01 181.13 27.62 ;
      RECT 180.39 21.01 181.13 21.21 ;
      RECT 180.39 18.71 180.59 21.21 ;
      RECT 179.09 37.61 179.69 37.81 ;
      RECT 179.49 27.02 179.69 37.81 ;
      RECT 179.49 27.02 180.73 27.22 ;
      RECT 180.53 21.41 180.73 27.22 ;
      RECT 179.99 21.41 180.73 21.61 ;
      RECT 179.99 12.98 180.19 21.61 ;
      RECT 180.13 21.81 180.33 23.85 ;
      RECT 179.59 21.81 180.33 22.01 ;
      RECT 179.59 20.73 179.79 22.01 ;
      RECT 179.49 38.01 179.69 65.05 ;
      RECT 179.49 38.01 180.09 38.21 ;
      RECT 179.89 30.13 180.09 38.21 ;
      RECT 176.29 67.59 180.09 68.59 ;
      RECT 177.99 26.07 178.39 68.59 ;
      RECT 177.49 26.07 178.39 28.61 ;
      RECT 177.49 26.07 178.89 28.6 ;
      RECT 176.83 26.07 179.55 26.27 ;
      RECT 179.35 24.87 179.55 26.27 ;
      RECT 176.83 24.87 177.03 26.27 ;
      RECT 176.83 24.87 179.55 25.07 ;
      RECT 177.49 14.44 178.89 25.07 ;
      RECT 177.99 6.24 178.39 25.07 ;
      RECT 177.69 6.24 179.19 6.84 ;
      RECT 179.09 38.01 179.29 65.45 ;
      RECT 178.69 38.01 179.29 38.21 ;
      RECT 178.69 30.13 178.89 38.21 ;
      RECT 178.39 510.34 179.19 510.94 ;
      RECT 177.19 510.34 177.99 510.94 ;
      RECT 177.19 510.34 179.19 510.74 ;
      RECT 176.69 37.61 177.29 37.81 ;
      RECT 176.69 27.02 176.89 37.81 ;
      RECT 175.65 27.02 176.89 27.22 ;
      RECT 175.65 21.41 175.85 27.22 ;
      RECT 175.65 21.41 176.39 21.61 ;
      RECT 176.19 19.42 176.39 21.61 ;
      RECT 176.19 19.42 176.99 19.62 ;
      RECT 176.79 13.78 176.99 19.62 ;
      RECT 176.79 13.78 177.79 13.98 ;
      RECT 177.59 8.94 177.79 13.98 ;
      RECT 177.09 38.01 177.29 65.45 ;
      RECT 177.09 38.01 177.69 38.21 ;
      RECT 177.49 30.13 177.69 38.21 ;
      RECT 175.59 27.82 175.99 68.59 ;
      RECT 173.89 65.96 177.69 66.96 ;
      RECT 174.85 27.82 175.99 28.22 ;
      RECT 174.85 7.54 175.05 28.22 ;
      RECT 174.85 16.1 175.59 20.81 ;
      RECT 174.45 14.76 175.19 16.84 ;
      RECT 174.85 7.54 175.59 15.5 ;
      RECT 175.29 6.24 176.09 8.24 ;
      RECT 175.29 6.24 176.29 6.84 ;
      RECT 177.19 8.94 177.39 13.58 ;
      RECT 176.92 8.94 177.39 9.14 ;
      RECT 176.69 38.01 176.89 65.05 ;
      RECT 176.29 38.01 176.89 38.21 ;
      RECT 176.29 30.13 176.49 38.21 ;
      RECT 176.05 21.81 176.25 23.85 ;
      RECT 176.05 21.81 176.79 22.01 ;
      RECT 176.59 20.73 176.79 22.01 ;
      RECT 176.19 27.42 176.39 28.57 ;
      RECT 175.25 27.42 176.39 27.62 ;
      RECT 175.25 21.01 175.45 27.62 ;
      RECT 175.25 21.01 175.99 21.21 ;
      RECT 175.79 15.7 175.99 21.21 ;
      RECT 175.39 15.7 175.99 15.9 ;
      RECT 174.69 38.01 174.89 65.05 ;
      RECT 174.69 38.01 175.29 38.21 ;
      RECT 175.09 30.13 175.29 38.21 ;
      RECT 171.49 67.59 175.29 68.59 ;
      RECT 173.19 6.24 173.59 68.59 ;
      RECT 174.29 37.61 174.89 37.81 ;
      RECT 174.69 28.55 174.89 37.81 ;
      RECT 171.89 37.61 172.49 37.81 ;
      RECT 171.89 28.55 172.09 37.81 ;
      RECT 174.29 28.55 174.49 37.41 ;
      RECT 172.29 28.55 172.49 37.41 ;
      RECT 172.29 28.55 174.49 28.95 ;
      RECT 171.89 28.55 174.89 28.75 ;
      RECT 172.99 6.24 173.79 6.84 ;
      RECT 173.79 9.82 173.99 15.58 ;
      RECT 173.79 9.82 174.49 10.02 ;
      RECT 174.29 7.14 174.49 10.02 ;
      RECT 174.29 38.01 174.49 65.45 ;
      RECT 173.89 38.01 174.49 38.21 ;
      RECT 173.89 30.13 174.09 38.21 ;
      RECT 174.04 25.29 174.24 28.35 ;
      RECT 174.04 25.29 174.45 25.49 ;
      RECT 174.25 21.25 174.45 25.49 ;
      RECT 173.59 510.34 174.39 510.94 ;
      RECT 172.39 510.34 173.19 510.94 ;
      RECT 172.39 510.34 174.39 510.74 ;
      RECT 172.79 9.82 172.99 15.58 ;
      RECT 172.29 9.82 172.99 10.02 ;
      RECT 172.29 7.14 172.49 10.02 ;
      RECT 172.29 38.01 172.49 65.45 ;
      RECT 172.29 38.01 172.89 38.21 ;
      RECT 172.69 30.13 172.89 38.21 ;
      RECT 170.79 27.82 171.19 68.59 ;
      RECT 169.09 65.96 172.89 66.96 ;
      RECT 170.79 27.82 171.93 28.22 ;
      RECT 171.73 7.54 171.93 28.22 ;
      RECT 171.19 16.1 171.93 20.81 ;
      RECT 171.59 14.76 172.33 16.84 ;
      RECT 171.19 7.54 171.93 15.5 ;
      RECT 170.69 6.24 171.49 8.24 ;
      RECT 170.49 6.24 171.49 6.84 ;
      RECT 172.54 25.29 172.74 28.35 ;
      RECT 172.33 25.29 172.74 25.49 ;
      RECT 172.33 21.25 172.53 25.49 ;
      RECT 171.89 38.01 172.09 65.05 ;
      RECT 171.49 38.01 172.09 38.21 ;
      RECT 171.49 30.13 171.69 38.21 ;
      RECT 170.39 27.42 170.59 28.57 ;
      RECT 170.39 27.42 171.53 27.62 ;
      RECT 171.33 21.01 171.53 27.62 ;
      RECT 170.79 21.01 171.53 21.21 ;
      RECT 170.79 15.7 170.99 21.21 ;
      RECT 170.79 15.7 171.39 15.9 ;
      RECT 169.49 37.61 170.09 37.81 ;
      RECT 169.89 27.02 170.09 37.81 ;
      RECT 169.89 27.02 171.13 27.22 ;
      RECT 170.93 21.41 171.13 27.22 ;
      RECT 170.39 21.41 171.13 21.61 ;
      RECT 170.39 19.42 170.59 21.61 ;
      RECT 169.79 19.42 170.59 19.62 ;
      RECT 169.79 13.78 169.99 19.62 ;
      RECT 168.99 13.78 169.99 13.98 ;
      RECT 168.99 8.94 169.19 13.98 ;
      RECT 170.53 21.81 170.73 23.85 ;
      RECT 169.99 21.81 170.73 22.01 ;
      RECT 169.99 20.73 170.19 22.01 ;
      RECT 169.89 38.01 170.09 65.05 ;
      RECT 169.89 38.01 170.49 38.21 ;
      RECT 170.29 30.13 170.49 38.21 ;
      RECT 166.69 67.59 170.49 68.59 ;
      RECT 168.39 26.07 168.79 68.59 ;
      RECT 168.39 26.07 169.29 28.61 ;
      RECT 167.89 26.07 169.29 28.6 ;
      RECT 167.23 26.07 169.95 26.27 ;
      RECT 169.75 24.87 169.95 26.27 ;
      RECT 167.23 24.87 167.43 26.27 ;
      RECT 167.23 24.87 169.95 25.07 ;
      RECT 167.89 14.44 169.29 25.07 ;
      RECT 168.39 6.24 168.79 25.07 ;
      RECT 167.59 6.24 169.09 6.84 ;
      RECT 169.39 8.94 169.59 13.58 ;
      RECT 169.39 8.94 169.86 9.14 ;
      RECT 169.49 38.01 169.69 65.45 ;
      RECT 169.09 38.01 169.69 38.21 ;
      RECT 169.09 30.13 169.29 38.21 ;
      RECT 168.79 510.34 169.59 510.94 ;
      RECT 167.59 510.34 168.39 510.94 ;
      RECT 167.59 510.34 169.59 510.74 ;
      RECT 167.49 38.01 167.69 65.45 ;
      RECT 167.49 38.01 168.09 38.21 ;
      RECT 167.89 30.13 168.09 38.21 ;
      RECT 165.99 27.82 166.39 68.59 ;
      RECT 164.29 65.96 168.09 66.96 ;
      RECT 165.25 27.82 166.39 28.22 ;
      RECT 165.25 7.54 165.45 28.22 ;
      RECT 165.25 7.54 165.99 20.81 ;
      RECT 165.59 6.24 166.39 8.24 ;
      RECT 165.19 6.24 167.16 6.84 ;
      RECT 167.09 37.61 167.69 37.81 ;
      RECT 167.09 27.02 167.29 37.81 ;
      RECT 166.05 27.02 167.29 27.22 ;
      RECT 166.05 21.41 166.25 27.22 ;
      RECT 166.05 21.41 166.79 21.61 ;
      RECT 166.59 12.98 166.79 21.61 ;
      RECT 167.09 38.01 167.29 65.05 ;
      RECT 166.69 38.01 167.29 38.21 ;
      RECT 166.69 30.13 166.89 38.21 ;
      RECT 166.45 21.81 166.65 23.85 ;
      RECT 166.45 21.81 167.19 22.01 ;
      RECT 166.99 20.73 167.19 22.01 ;
      RECT 166.59 27.42 166.79 28.57 ;
      RECT 165.65 27.42 166.79 27.62 ;
      RECT 165.65 21.01 165.85 27.62 ;
      RECT 165.65 21.01 166.39 21.21 ;
      RECT 166.19 18.71 166.39 21.21 ;
      RECT 165.09 38.01 165.29 65.05 ;
      RECT 165.09 38.01 165.69 38.21 ;
      RECT 165.49 30.13 165.69 38.21 ;
      RECT 161.89 67.59 165.69 68.59 ;
      RECT 163.59 6.24 163.99 68.59 ;
      RECT 164.69 37.61 165.29 37.81 ;
      RECT 165.09 28.55 165.29 37.81 ;
      RECT 162.29 37.61 162.89 37.81 ;
      RECT 162.29 28.55 162.49 37.81 ;
      RECT 164.69 28.55 164.89 37.41 ;
      RECT 162.69 28.55 162.89 37.41 ;
      RECT 163.59 28.55 164.89 28.95 ;
      RECT 162.29 28.55 165.29 28.75 ;
      RECT 162.89 28.15 163.99 28.75 ;
      RECT 163.59 9.34 164.39 9.54 ;
      RECT 162.79 6.24 164.79 6.84 ;
      RECT 164.69 38.01 164.89 65.45 ;
      RECT 164.29 38.01 164.89 38.21 ;
      RECT 164.29 30.13 164.49 38.21 ;
      RECT 164.44 25.29 164.64 28.35 ;
      RECT 164.44 25.29 164.85 25.49 ;
      RECT 164.65 21.25 164.85 25.49 ;
      RECT 163.99 510.34 164.79 510.94 ;
      RECT 162.79 510.34 163.59 510.94 ;
      RECT 162.79 510.34 164.79 510.74 ;
      RECT 162.69 38.01 162.89 65.45 ;
      RECT 162.69 38.01 163.29 38.21 ;
      RECT 163.09 30.13 163.29 38.21 ;
      RECT 161.19 27.82 161.59 68.59 ;
      RECT 159.49 65.96 163.29 66.96 ;
      RECT 161.59 6.24 162.33 28.22 ;
      RECT 160.39 6.24 162.33 18.31 ;
      RECT 160.39 6.24 162.37 7.44 ;
      RECT 162.29 38.01 162.49 65.05 ;
      RECT 161.89 38.01 162.49 38.21 ;
      RECT 161.89 30.13 162.09 38.21 ;
      RECT 160.29 38.01 160.49 65.05 ;
      RECT 160.29 38.01 160.89 38.21 ;
      RECT 160.69 30.13 160.89 38.21 ;
      RECT 157.09 67.59 160.89 68.59 ;
      RECT 158.79 28.15 159.19 68.59 ;
      RECT 159.89 37.61 160.49 37.81 ;
      RECT 160.29 28.75 160.49 37.81 ;
      RECT 159.89 28.15 160.09 37.41 ;
      RECT 159.89 28.75 160.49 28.95 ;
      RECT 159.89 38.01 160.09 65.45 ;
      RECT 159.49 38.01 160.09 38.21 ;
      RECT 159.49 30.13 159.69 38.21 ;
      RECT 159.19 510.34 159.99 510.94 ;
      RECT 157.99 510.34 158.79 510.94 ;
      RECT 157.99 510.34 159.99 510.74 ;
      RECT 158.29 6.24 159.69 25.07 ;
      RECT 157.99 6.24 159.97 7.44 ;
      RECT 157.89 38.01 158.09 65.45 ;
      RECT 157.89 38.01 158.49 38.21 ;
      RECT 158.29 30.13 158.49 38.21 ;
      RECT 156.39 27.82 156.79 68.59 ;
      RECT 154.69 65.96 158.49 66.96 ;
      RECT 155.65 6.24 156.39 28.22 ;
      RECT 155.65 6.24 157.57 18.31 ;
      RECT 155.59 6.24 157.57 7.44 ;
      RECT 157.49 37.61 158.09 37.81 ;
      RECT 157.49 28.75 157.69 37.81 ;
      RECT 157.89 28.15 158.09 37.41 ;
      RECT 157.49 28.75 158.09 28.95 ;
      RECT 157.49 38.01 157.69 65.05 ;
      RECT 157.09 38.01 157.69 38.21 ;
      RECT 157.09 30.13 157.29 38.21 ;
      RECT 155.49 38.01 155.69 65.05 ;
      RECT 155.49 38.01 156.09 38.21 ;
      RECT 155.89 30.13 156.09 38.21 ;
      RECT 153.99 67.59 156.09 68.59 ;
      RECT 153.99 6.24 154.39 68.59 ;
      RECT 155.09 37.61 155.69 37.81 ;
      RECT 155.49 28.55 155.69 37.81 ;
      RECT 155.09 28.55 155.29 37.41 ;
      RECT 153.99 28.55 155.69 28.75 ;
      RECT 153.99 28.15 155.09 28.75 ;
      RECT 153.89 6.24 155.19 6.84 ;
      RECT 155.09 38.01 155.29 65.45 ;
      RECT 154.69 38.01 155.29 38.21 ;
      RECT 154.69 30.13 154.89 38.21 ;
      RECT 154.39 510.34 155.19 510.94 ;
      RECT 153.19 510.34 153.99 510.94 ;
      RECT 153.19 510.34 155.19 510.74 ;
      RECT 152.89 23.14 153.09 43.05 ;
      RECT 152.89 23.14 153.49 23.34 ;
      RECT 153.29 7.14 153.49 23.34 ;
      RECT 152.69 67.98 152.89 68.66 ;
      RECT 152.69 67.98 153.49 68.18 ;
      RECT 153.29 23.74 153.49 68.18 ;
      RECT 151.69 6.24 151.89 27.71 ;
      RECT 151.29 6.24 151.89 6.84 ;
      RECT 151.59 31.23 151.79 51.87 ;
      RECT 150.89 31.23 151.79 31.43 ;
      RECT 150.89 25.43 151.09 31.43 ;
      RECT 149.93 32.39 150.49 69.03 ;
      RECT 150.29 6.24 150.69 66.83 ;
      RECT 150.29 6.24 150.89 8.59 ;
      RECT 146.09 32.39 147.41 510.94 ;
      RECT 146.55 6.24 146.95 510.94 ;
      RECT 146.09 6.24 147.41 6.84 ;
      RECT 144.17 32.39 145.49 510.94 ;
      RECT 144.63 8.19 145.03 510.94 ;
      RECT 145.01 6.24 145.61 8.59 ;
      RECT 142.25 32.39 143.57 510.94 ;
      RECT 142.71 6.24 143.11 510.94 ;
      RECT 142.62 6.24 143.57 8.56 ;
      RECT 141.99 6.24 142.22 29.57 ;
      RECT 141.62 6.24 142.22 6.84 ;
      RECT 138.41 69.46 141.65 510.94 ;
      RECT 140.79 32.39 141.65 510.94 ;
      RECT 138.81 66.63 141.65 510.94 ;
      RECT 138.81 15.28 140.01 510.94 ;
      RECT 138.83 6.24 140.01 510.94 ;
      RECT 140.79 8.19 141.19 510.94 ;
      RECT 138.83 6.24 140.81 11.84 ;
      RECT 138.83 6.24 140.83 6.84 ;
      RECT 135.01 69.56 137.81 510.94 ;
      RECT 135.41 15.28 137.41 510.94 ;
      RECT 135.43 6.24 137.39 510.94 ;
      RECT 134.81 48.74 135.01 49.84 ;
      RECT 134.61 16.13 134.81 48.94 ;
      RECT 134.61 50.04 134.81 65.83 ;
      RECT 134.41 49.14 134.61 50.24 ;
      RECT 131.61 69.46 134.41 510.94 ;
      RECT 132.01 39.44 134.01 510.94 ;
      RECT 132.81 6.24 133.21 510.94 ;
      RECT 132.01 15.28 134.01 32.15 ;
      RECT 132.03 6.24 133.99 32.15 ;
      RECT 132.12 34.93 132.32 38.18 ;
      RECT 131.61 34.93 132.32 35.13 ;
      RECT 131.61 12.32 131.81 35.13 ;
      RECT 131.41 47.54 131.61 48.64 ;
      RECT 131.21 16.13 131.41 47.74 ;
      RECT 131.21 48.84 131.41 65.83 ;
      RECT 131.01 47.94 131.21 49.04 ;
      RECT 128.21 69.46 131.01 510.94 ;
      RECT 128.61 39.44 130.61 510.94 ;
      RECT 129.41 6.24 129.81 510.94 ;
      RECT 128.61 15.28 130.61 32.15 ;
      RECT 128.63 6.24 130.59 32.15 ;
      RECT 128.01 46.34 128.21 47.44 ;
      RECT 127.81 16.13 128.01 46.54 ;
      RECT 127.81 47.64 128.01 65.83 ;
      RECT 127.61 46.74 127.81 47.84 ;
      RECT 124.81 69.56 127.61 510.94 ;
      RECT 125.21 39.44 127.21 510.94 ;
      RECT 126.01 6.24 126.41 510.94 ;
      RECT 125.21 15.28 127.21 32.15 ;
      RECT 125.21 6.24 127.19 32.15 ;
      RECT 124.61 45.14 124.81 46.24 ;
      RECT 124.41 16.13 124.61 45.34 ;
      RECT 124.41 46.44 124.61 65.83 ;
      RECT 124.21 45.54 124.41 46.64 ;
      RECT 122.61 6.24 123.01 66.63 ;
      RECT 122.61 6.24 123.81 65.33 ;
      RECT 122.31 41.29 123.81 54.42 ;
      RECT 121.83 6.24 123.81 32.15 ;
      RECT 121.23 66.03 121.73 66.43 ;
      RECT 121.43 54.14 121.73 66.43 ;
      RECT 121.01 54.14 121.73 54.44 ;
      RECT 121.01 44.24 121.31 54.44 ;
      RECT 121.01 16.13 121.21 54.44 ;
      RECT 120.46 65.53 120.94 66.43 ;
      RECT 120.46 65.53 121.21 65.83 ;
      RECT 121.01 61.91 121.21 65.83 ;
      RECT 118.01 505.69 120.81 510.94 ;
      RECT 118.91 39.44 119.91 510.94 ;
      RECT 119.21 6.24 119.61 510.94 ;
      RECT 118.43 6.24 120.39 32.15 ;
      RECT 118.52 34.93 118.72 38.18 ;
      RECT 118.01 34.93 118.72 35.13 ;
      RECT 118.01 12.32 118.21 35.13 ;
      RECT 117.84 66.04 118.49 66.43 ;
      RECT 118.19 61.1 118.49 66.43 ;
      RECT 117.52 61.1 118.49 61.4 ;
      RECT 117.52 44.24 117.82 61.4 ;
      RECT 117.61 16.13 117.81 61.4 ;
      RECT 117.06 65.53 117.54 66.43 ;
      RECT 117.06 65.53 117.81 65.83 ;
      RECT 117.61 61.91 117.81 65.83 ;
      RECT 114.61 505.69 117.41 510.94 ;
      RECT 115.51 39.44 116.51 510.94 ;
      RECT 115.81 6.24 116.21 510.94 ;
      RECT 115.03 6.24 116.99 32.15 ;
      RECT 114.43 66.03 114.93 66.43 ;
      RECT 114.63 54.14 114.93 66.43 ;
      RECT 114.21 54.14 114.93 54.44 ;
      RECT 114.21 44.24 114.51 54.44 ;
      RECT 114.21 16.13 114.41 54.44 ;
      RECT 113.66 65.53 114.14 66.43 ;
      RECT 113.66 65.53 114.41 65.83 ;
      RECT 114.21 61.91 114.41 65.83 ;
      RECT 111.21 505.69 114.01 510.94 ;
      RECT 112.11 39.44 113.11 510.94 ;
      RECT 112.41 6.24 112.81 510.94 ;
      RECT 111.61 6.24 113.59 32.15 ;
      RECT 111.03 66.03 111.69 66.43 ;
      RECT 111.39 61.1 111.69 66.43 ;
      RECT 110.72 61.1 111.69 61.4 ;
      RECT 110.72 44.24 111.02 61.4 ;
      RECT 110.81 16.13 111.01 61.4 ;
      RECT 110.26 65.53 110.74 66.43 ;
      RECT 110.26 65.53 111.01 65.83 ;
      RECT 110.81 61.91 111.01 65.83 ;
      RECT 109.01 6.24 109.41 66.63 ;
      RECT 108.71 41.29 109.71 54.42 ;
      RECT 109.01 39.44 109.71 54.42 ;
      RECT 108.23 6.24 110.21 32.15 ;
      RECT 7.2 70.16 110.06 70.66 ;
      RECT 109.46 69.86 110.06 70.66 ;
      RECT 109.46 71.86 110.06 72.67 ;
      RECT 7.2 71.86 110.06 72.36 ;
      RECT 7.2 73.56 110.06 74.06 ;
      RECT 109.46 73.25 110.06 74.06 ;
      RECT 109.46 75.26 110.06 76.06 ;
      RECT 7.2 75.26 110.06 75.76 ;
      RECT 7.2 76.96 110.06 77.46 ;
      RECT 109.46 76.66 110.06 77.46 ;
      RECT 109.46 78.66 110.06 79.47 ;
      RECT 7.2 78.66 110.06 79.16 ;
      RECT 7.2 80.36 110.06 80.86 ;
      RECT 109.46 80.05 110.06 80.86 ;
      RECT 109.46 82.06 110.06 82.86 ;
      RECT 7.2 82.06 110.06 82.56 ;
      RECT 7.2 83.76 110.06 84.26 ;
      RECT 109.46 83.46 110.06 84.26 ;
      RECT 109.46 85.46 110.06 86.27 ;
      RECT 7.2 85.46 110.06 85.96 ;
      RECT 7.2 87.16 110.06 87.66 ;
      RECT 109.46 86.85 110.06 87.66 ;
      RECT 109.46 88.86 110.06 89.66 ;
      RECT 7.2 88.86 110.06 89.36 ;
      RECT 7.2 90.56 110.06 91.06 ;
      RECT 109.46 90.26 110.06 91.06 ;
      RECT 109.46 92.26 110.06 93.07 ;
      RECT 7.2 92.26 110.06 92.76 ;
      RECT 7.2 93.96 110.06 94.46 ;
      RECT 109.46 93.65 110.06 94.46 ;
      RECT 109.46 95.66 110.06 96.46 ;
      RECT 7.2 95.66 110.06 96.16 ;
      RECT 7.2 97.36 110.06 97.86 ;
      RECT 109.46 97.06 110.06 97.86 ;
      RECT 109.46 99.06 110.06 99.87 ;
      RECT 7.2 99.06 110.06 99.56 ;
      RECT 7.2 100.76 110.06 101.26 ;
      RECT 109.46 100.45 110.06 101.26 ;
      RECT 109.46 102.46 110.06 103.26 ;
      RECT 7.2 102.46 110.06 102.96 ;
      RECT 7.2 104.16 110.06 104.66 ;
      RECT 109.46 103.86 110.06 104.66 ;
      RECT 109.46 105.86 110.06 106.67 ;
      RECT 7.2 105.86 110.06 106.36 ;
      RECT 7.2 107.56 110.06 108.06 ;
      RECT 109.46 107.25 110.06 108.06 ;
      RECT 109.46 109.26 110.06 110.06 ;
      RECT 7.2 109.26 110.06 109.76 ;
      RECT 7.2 110.96 110.06 111.46 ;
      RECT 109.46 110.66 110.06 111.46 ;
      RECT 109.46 112.66 110.06 113.47 ;
      RECT 7.2 112.66 110.06 113.16 ;
      RECT 7.2 114.36 110.06 114.86 ;
      RECT 109.46 114.05 110.06 114.86 ;
      RECT 109.46 116.06 110.06 116.86 ;
      RECT 7.2 116.06 110.06 116.56 ;
      RECT 7.2 117.76 110.06 118.26 ;
      RECT 109.46 117.46 110.06 118.26 ;
      RECT 109.46 119.46 110.06 120.27 ;
      RECT 7.2 119.46 110.06 119.96 ;
      RECT 7.2 121.16 110.06 121.66 ;
      RECT 109.46 120.85 110.06 121.66 ;
      RECT 109.46 122.86 110.06 123.66 ;
      RECT 7.2 122.86 110.06 123.36 ;
      RECT 7.2 124.56 110.06 125.06 ;
      RECT 109.46 124.26 110.06 125.06 ;
      RECT 109.46 126.26 110.06 127.07 ;
      RECT 7.2 126.26 110.06 126.76 ;
      RECT 7.2 127.96 110.06 128.46 ;
      RECT 109.46 127.65 110.06 128.46 ;
      RECT 109.46 129.66 110.06 130.46 ;
      RECT 7.2 129.66 110.06 130.16 ;
      RECT 7.2 131.36 110.06 131.86 ;
      RECT 109.46 131.06 110.06 131.86 ;
      RECT 109.46 133.06 110.06 133.87 ;
      RECT 7.2 133.06 110.06 133.56 ;
      RECT 7.2 134.76 110.06 135.26 ;
      RECT 109.46 134.45 110.06 135.26 ;
      RECT 109.46 136.46 110.06 137.26 ;
      RECT 7.2 136.46 110.06 136.96 ;
      RECT 7.2 138.16 110.06 138.66 ;
      RECT 109.46 137.86 110.06 138.66 ;
      RECT 109.46 139.86 110.06 140.67 ;
      RECT 7.2 139.86 110.06 140.36 ;
      RECT 7.2 141.56 110.06 142.06 ;
      RECT 109.46 141.25 110.06 142.06 ;
      RECT 109.46 143.26 110.06 144.06 ;
      RECT 7.2 143.26 110.06 143.76 ;
      RECT 7.2 144.96 110.06 145.46 ;
      RECT 109.46 144.66 110.06 145.46 ;
      RECT 109.46 146.66 110.06 147.47 ;
      RECT 7.2 146.66 110.06 147.16 ;
      RECT 7.2 148.36 110.06 148.86 ;
      RECT 109.46 148.05 110.06 148.86 ;
      RECT 109.46 150.06 110.06 150.86 ;
      RECT 7.2 150.06 110.06 150.56 ;
      RECT 7.2 151.76 110.06 152.26 ;
      RECT 109.46 151.46 110.06 152.26 ;
      RECT 109.46 153.46 110.06 154.27 ;
      RECT 7.2 153.46 110.06 153.96 ;
      RECT 7.2 155.16 110.06 155.66 ;
      RECT 109.46 154.85 110.06 155.66 ;
      RECT 109.46 156.86 110.06 157.66 ;
      RECT 7.2 156.86 110.06 157.36 ;
      RECT 7.2 158.56 110.06 159.06 ;
      RECT 109.46 158.26 110.06 159.06 ;
      RECT 109.46 160.26 110.06 161.07 ;
      RECT 7.2 160.26 110.06 160.76 ;
      RECT 7.2 161.96 110.06 162.46 ;
      RECT 109.46 161.65 110.06 162.46 ;
      RECT 109.46 163.66 110.06 164.46 ;
      RECT 7.2 163.66 110.06 164.16 ;
      RECT 7.2 165.36 110.06 165.86 ;
      RECT 109.46 165.06 110.06 165.86 ;
      RECT 109.46 167.06 110.06 167.87 ;
      RECT 7.2 167.06 110.06 167.56 ;
      RECT 7.2 168.76 110.06 169.26 ;
      RECT 109.46 168.45 110.06 169.26 ;
      RECT 109.46 170.46 110.06 171.26 ;
      RECT 7.2 170.46 110.06 170.96 ;
      RECT 7.2 172.16 110.06 172.66 ;
      RECT 109.46 171.86 110.06 172.66 ;
      RECT 109.46 173.86 110.06 174.67 ;
      RECT 7.2 173.86 110.06 174.36 ;
      RECT 7.2 175.56 110.06 176.06 ;
      RECT 109.46 175.25 110.06 176.06 ;
      RECT 109.46 177.26 110.06 178.06 ;
      RECT 7.2 177.26 110.06 177.76 ;
      RECT 7.2 178.96 110.06 179.46 ;
      RECT 109.46 178.66 110.06 179.46 ;
      RECT 109.46 180.66 110.06 181.47 ;
      RECT 7.2 180.66 110.06 181.16 ;
      RECT 7.2 182.36 110.06 182.86 ;
      RECT 109.46 182.05 110.06 182.86 ;
      RECT 109.46 184.06 110.06 184.86 ;
      RECT 7.2 184.06 110.06 184.56 ;
      RECT 7.2 185.76 110.06 186.26 ;
      RECT 109.46 185.46 110.06 186.26 ;
      RECT 109.46 187.46 110.06 188.27 ;
      RECT 7.2 187.46 110.06 187.96 ;
      RECT 7.2 189.16 110.06 189.66 ;
      RECT 109.46 188.85 110.06 189.66 ;
      RECT 109.46 190.86 110.06 191.66 ;
      RECT 7.2 190.86 110.06 191.36 ;
      RECT 7.2 192.56 110.06 193.06 ;
      RECT 109.46 192.26 110.06 193.06 ;
      RECT 109.46 194.26 110.06 195.07 ;
      RECT 7.2 194.26 110.06 194.76 ;
      RECT 7.2 195.96 110.06 196.46 ;
      RECT 109.46 195.65 110.06 196.46 ;
      RECT 109.46 197.66 110.06 198.46 ;
      RECT 7.2 197.66 110.06 198.16 ;
      RECT 7.2 199.36 110.06 199.86 ;
      RECT 109.46 199.06 110.06 199.86 ;
      RECT 109.46 201.06 110.06 201.87 ;
      RECT 7.2 201.06 110.06 201.56 ;
      RECT 7.2 202.76 110.06 203.26 ;
      RECT 109.46 202.45 110.06 203.26 ;
      RECT 109.46 204.46 110.06 205.26 ;
      RECT 7.2 204.46 110.06 204.96 ;
      RECT 7.2 206.16 110.06 206.66 ;
      RECT 109.46 205.86 110.06 206.66 ;
      RECT 109.46 207.86 110.06 208.67 ;
      RECT 7.2 207.86 110.06 208.36 ;
      RECT 7.2 209.56 110.06 210.06 ;
      RECT 109.46 209.25 110.06 210.06 ;
      RECT 109.46 211.26 110.06 212.06 ;
      RECT 7.2 211.26 110.06 211.76 ;
      RECT 7.2 212.96 110.06 213.46 ;
      RECT 109.46 212.66 110.06 213.46 ;
      RECT 109.46 214.66 110.06 215.47 ;
      RECT 7.2 214.66 110.06 215.16 ;
      RECT 7.2 216.36 110.06 216.86 ;
      RECT 109.46 216.05 110.06 216.86 ;
      RECT 109.46 218.06 110.06 218.86 ;
      RECT 7.2 218.06 110.06 218.56 ;
      RECT 7.2 219.76 110.06 220.26 ;
      RECT 109.46 219.46 110.06 220.26 ;
      RECT 109.46 221.46 110.06 222.27 ;
      RECT 7.2 221.46 110.06 221.96 ;
      RECT 7.2 223.16 110.06 223.66 ;
      RECT 109.46 222.85 110.06 223.66 ;
      RECT 109.46 224.86 110.06 225.66 ;
      RECT 7.2 224.86 110.06 225.36 ;
      RECT 7.2 226.56 110.06 227.06 ;
      RECT 109.46 226.26 110.06 227.06 ;
      RECT 109.46 228.26 110.06 229.07 ;
      RECT 7.2 228.26 110.06 228.76 ;
      RECT 7.2 229.96 110.06 230.46 ;
      RECT 109.46 229.65 110.06 230.46 ;
      RECT 109.46 231.66 110.06 232.46 ;
      RECT 7.2 231.66 110.06 232.16 ;
      RECT 7.2 233.36 110.06 233.86 ;
      RECT 109.46 233.06 110.06 233.86 ;
      RECT 109.46 235.06 110.06 235.87 ;
      RECT 7.2 235.06 110.06 235.56 ;
      RECT 7.2 236.76 110.06 237.26 ;
      RECT 109.46 236.45 110.06 237.26 ;
      RECT 109.46 238.46 110.06 239.26 ;
      RECT 7.2 238.46 110.06 238.96 ;
      RECT 7.2 240.16 110.06 240.66 ;
      RECT 109.46 239.86 110.06 240.66 ;
      RECT 109.46 241.86 110.06 242.67 ;
      RECT 7.2 241.86 110.06 242.36 ;
      RECT 7.2 243.56 110.06 244.06 ;
      RECT 109.46 243.25 110.06 244.06 ;
      RECT 109.46 245.26 110.06 246.06 ;
      RECT 7.2 245.26 110.06 245.76 ;
      RECT 7.2 246.96 110.06 247.46 ;
      RECT 109.46 246.66 110.06 247.46 ;
      RECT 109.46 248.66 110.06 249.47 ;
      RECT 7.2 248.66 110.06 249.16 ;
      RECT 7.2 250.36 110.06 250.86 ;
      RECT 109.46 250.05 110.06 250.86 ;
      RECT 109.46 252.06 110.06 252.86 ;
      RECT 7.2 252.06 110.06 252.56 ;
      RECT 7.2 253.76 110.06 254.26 ;
      RECT 109.46 253.46 110.06 254.26 ;
      RECT 109.46 255.46 110.06 256.27 ;
      RECT 7.2 255.46 110.06 255.96 ;
      RECT 7.2 257.16 110.06 257.66 ;
      RECT 109.46 256.85 110.06 257.66 ;
      RECT 109.46 258.86 110.06 259.66 ;
      RECT 7.2 258.86 110.06 259.36 ;
      RECT 7.2 260.56 110.06 261.06 ;
      RECT 109.46 260.26 110.06 261.06 ;
      RECT 109.46 262.26 110.06 263.07 ;
      RECT 7.2 262.26 110.06 262.76 ;
      RECT 7.2 263.96 110.06 264.46 ;
      RECT 109.46 263.65 110.06 264.46 ;
      RECT 109.46 265.66 110.06 266.46 ;
      RECT 7.2 265.66 110.06 266.16 ;
      RECT 7.2 267.36 110.06 267.86 ;
      RECT 109.46 267.06 110.06 267.86 ;
      RECT 109.46 269.06 110.06 269.87 ;
      RECT 7.2 269.06 110.06 269.56 ;
      RECT 7.2 270.76 110.06 271.26 ;
      RECT 109.46 270.45 110.06 271.26 ;
      RECT 109.46 272.46 110.06 273.26 ;
      RECT 7.2 272.46 110.06 272.96 ;
      RECT 7.2 274.16 110.06 274.66 ;
      RECT 109.46 273.86 110.06 274.66 ;
      RECT 109.46 275.86 110.06 276.67 ;
      RECT 7.2 275.86 110.06 276.36 ;
      RECT 7.2 277.56 110.06 278.06 ;
      RECT 109.46 277.25 110.06 278.06 ;
      RECT 109.46 279.26 110.06 280.06 ;
      RECT 7.2 279.26 110.06 279.76 ;
      RECT 7.2 280.96 110.06 281.46 ;
      RECT 109.46 280.66 110.06 281.46 ;
      RECT 109.46 282.66 110.06 283.47 ;
      RECT 7.2 282.66 110.06 283.16 ;
      RECT 7.2 284.36 110.06 284.86 ;
      RECT 109.46 284.05 110.06 284.86 ;
      RECT 109.46 286.06 110.06 286.86 ;
      RECT 7.2 286.06 110.06 286.56 ;
      RECT 7.2 287.76 110.06 288.26 ;
      RECT 109.46 287.46 110.06 288.26 ;
      RECT 109.46 289.46 110.06 290.27 ;
      RECT 7.2 289.46 110.06 289.96 ;
      RECT 7.2 291.16 110.06 291.66 ;
      RECT 109.46 290.85 110.06 291.66 ;
      RECT 109.46 292.86 110.06 293.66 ;
      RECT 7.2 292.86 110.06 293.36 ;
      RECT 7.2 294.56 110.06 295.06 ;
      RECT 109.46 294.26 110.06 295.06 ;
      RECT 109.46 296.26 110.06 297.07 ;
      RECT 7.2 296.26 110.06 296.76 ;
      RECT 7.2 297.96 110.06 298.46 ;
      RECT 109.46 297.65 110.06 298.46 ;
      RECT 109.46 299.66 110.06 300.46 ;
      RECT 7.2 299.66 110.06 300.16 ;
      RECT 7.2 301.36 110.06 301.86 ;
      RECT 109.46 301.06 110.06 301.86 ;
      RECT 109.46 303.06 110.06 303.87 ;
      RECT 7.2 303.06 110.06 303.56 ;
      RECT 7.2 304.76 110.06 305.26 ;
      RECT 109.46 304.45 110.06 305.26 ;
      RECT 109.46 306.46 110.06 307.26 ;
      RECT 7.2 306.46 110.06 306.96 ;
      RECT 7.2 308.16 110.06 308.66 ;
      RECT 109.46 307.86 110.06 308.66 ;
      RECT 109.46 309.86 110.06 310.67 ;
      RECT 7.2 309.86 110.06 310.36 ;
      RECT 7.2 311.56 110.06 312.06 ;
      RECT 109.46 311.25 110.06 312.06 ;
      RECT 109.46 313.26 110.06 314.06 ;
      RECT 7.2 313.26 110.06 313.76 ;
      RECT 7.2 314.96 110.06 315.46 ;
      RECT 109.46 314.66 110.06 315.46 ;
      RECT 109.46 316.66 110.06 317.47 ;
      RECT 7.2 316.66 110.06 317.16 ;
      RECT 7.2 318.36 110.06 318.86 ;
      RECT 109.46 318.05 110.06 318.86 ;
      RECT 109.46 320.06 110.06 320.86 ;
      RECT 7.2 320.06 110.06 320.56 ;
      RECT 7.2 321.76 110.06 322.26 ;
      RECT 109.46 321.46 110.06 322.26 ;
      RECT 109.46 323.46 110.06 324.27 ;
      RECT 7.2 323.46 110.06 323.96 ;
      RECT 7.2 325.16 110.06 325.66 ;
      RECT 109.46 324.85 110.06 325.66 ;
      RECT 109.46 326.86 110.06 327.66 ;
      RECT 7.2 326.86 110.06 327.36 ;
      RECT 7.2 328.56 110.06 329.06 ;
      RECT 109.46 328.26 110.06 329.06 ;
      RECT 109.46 330.26 110.06 331.07 ;
      RECT 7.2 330.26 110.06 330.76 ;
      RECT 7.2 331.96 110.06 332.46 ;
      RECT 109.46 331.65 110.06 332.46 ;
      RECT 109.46 333.66 110.06 334.46 ;
      RECT 7.2 333.66 110.06 334.16 ;
      RECT 7.2 335.36 110.06 335.86 ;
      RECT 109.46 335.06 110.06 335.86 ;
      RECT 109.46 337.06 110.06 337.87 ;
      RECT 7.2 337.06 110.06 337.56 ;
      RECT 7.2 338.76 110.06 339.26 ;
      RECT 109.46 338.45 110.06 339.26 ;
      RECT 109.46 340.46 110.06 341.26 ;
      RECT 7.2 340.46 110.06 340.96 ;
      RECT 7.2 342.16 110.06 342.66 ;
      RECT 109.46 341.86 110.06 342.66 ;
      RECT 109.46 343.86 110.06 344.67 ;
      RECT 7.2 343.86 110.06 344.36 ;
      RECT 7.2 345.56 110.06 346.06 ;
      RECT 109.46 345.25 110.06 346.06 ;
      RECT 109.46 347.26 110.06 348.06 ;
      RECT 7.2 347.26 110.06 347.76 ;
      RECT 7.2 348.96 110.06 349.46 ;
      RECT 109.46 348.66 110.06 349.46 ;
      RECT 109.46 350.66 110.06 351.47 ;
      RECT 7.2 350.66 110.06 351.16 ;
      RECT 7.2 352.36 110.06 352.86 ;
      RECT 109.46 352.05 110.06 352.86 ;
      RECT 109.46 354.06 110.06 354.86 ;
      RECT 7.2 354.06 110.06 354.56 ;
      RECT 7.2 355.76 110.06 356.26 ;
      RECT 109.46 355.46 110.06 356.26 ;
      RECT 109.46 357.46 110.06 358.27 ;
      RECT 7.2 357.46 110.06 357.96 ;
      RECT 7.2 359.16 110.06 359.66 ;
      RECT 109.46 358.85 110.06 359.66 ;
      RECT 109.46 360.86 110.06 361.66 ;
      RECT 7.2 360.86 110.06 361.36 ;
      RECT 7.2 362.56 110.06 363.06 ;
      RECT 109.46 362.26 110.06 363.06 ;
      RECT 109.46 364.26 110.06 365.07 ;
      RECT 7.2 364.26 110.06 364.76 ;
      RECT 7.2 365.96 110.06 366.46 ;
      RECT 109.46 365.65 110.06 366.46 ;
      RECT 109.46 367.66 110.06 368.46 ;
      RECT 7.2 367.66 110.06 368.16 ;
      RECT 7.2 369.36 110.06 369.86 ;
      RECT 109.46 369.06 110.06 369.86 ;
      RECT 109.46 371.06 110.06 371.87 ;
      RECT 7.2 371.06 110.06 371.56 ;
      RECT 7.2 372.76 110.06 373.26 ;
      RECT 109.46 372.45 110.06 373.26 ;
      RECT 109.46 374.46 110.06 375.26 ;
      RECT 7.2 374.46 110.06 374.96 ;
      RECT 7.2 376.16 110.06 376.66 ;
      RECT 109.46 375.86 110.06 376.66 ;
      RECT 109.46 377.86 110.06 378.67 ;
      RECT 7.2 377.86 110.06 378.36 ;
      RECT 7.2 379.56 110.06 380.06 ;
      RECT 109.46 379.25 110.06 380.06 ;
      RECT 109.46 381.26 110.06 382.06 ;
      RECT 7.2 381.26 110.06 381.76 ;
      RECT 7.2 382.96 110.06 383.46 ;
      RECT 109.46 382.66 110.06 383.46 ;
      RECT 109.46 384.66 110.06 385.47 ;
      RECT 7.2 384.66 110.06 385.16 ;
      RECT 7.2 386.36 110.06 386.86 ;
      RECT 109.46 386.05 110.06 386.86 ;
      RECT 109.46 388.06 110.06 388.86 ;
      RECT 7.2 388.06 110.06 388.56 ;
      RECT 7.2 389.76 110.06 390.26 ;
      RECT 109.46 389.46 110.06 390.26 ;
      RECT 109.46 391.46 110.06 392.27 ;
      RECT 7.2 391.46 110.06 391.96 ;
      RECT 7.2 393.16 110.06 393.66 ;
      RECT 109.46 392.85 110.06 393.66 ;
      RECT 109.46 394.86 110.06 395.66 ;
      RECT 7.2 394.86 110.06 395.36 ;
      RECT 7.2 396.56 110.06 397.06 ;
      RECT 109.46 396.26 110.06 397.06 ;
      RECT 109.46 398.26 110.06 399.07 ;
      RECT 7.2 398.26 110.06 398.76 ;
      RECT 7.2 399.96 110.06 400.46 ;
      RECT 109.46 399.65 110.06 400.46 ;
      RECT 109.46 401.66 110.06 402.46 ;
      RECT 7.2 401.66 110.06 402.16 ;
      RECT 7.2 403.36 110.06 403.86 ;
      RECT 109.46 403.06 110.06 403.86 ;
      RECT 109.46 405.06 110.06 405.87 ;
      RECT 7.2 405.06 110.06 405.56 ;
      RECT 7.2 406.76 110.06 407.26 ;
      RECT 109.46 406.45 110.06 407.26 ;
      RECT 109.46 408.46 110.06 409.26 ;
      RECT 7.2 408.46 110.06 408.96 ;
      RECT 7.2 410.16 110.06 410.66 ;
      RECT 109.46 409.86 110.06 410.66 ;
      RECT 109.46 411.86 110.06 412.67 ;
      RECT 7.2 411.86 110.06 412.36 ;
      RECT 7.2 413.56 110.06 414.06 ;
      RECT 109.46 413.25 110.06 414.06 ;
      RECT 109.46 415.26 110.06 416.06 ;
      RECT 7.2 415.26 110.06 415.76 ;
      RECT 7.2 416.96 110.06 417.46 ;
      RECT 109.46 416.66 110.06 417.46 ;
      RECT 109.46 418.66 110.06 419.47 ;
      RECT 7.2 418.66 110.06 419.16 ;
      RECT 7.2 420.36 110.06 420.86 ;
      RECT 109.46 420.05 110.06 420.86 ;
      RECT 109.46 422.06 110.06 422.86 ;
      RECT 7.2 422.06 110.06 422.56 ;
      RECT 7.2 423.76 110.06 424.26 ;
      RECT 109.46 423.46 110.06 424.26 ;
      RECT 109.46 425.46 110.06 426.27 ;
      RECT 7.2 425.46 110.06 425.96 ;
      RECT 7.2 427.16 110.06 427.66 ;
      RECT 109.46 426.85 110.06 427.66 ;
      RECT 109.46 428.86 110.06 429.66 ;
      RECT 7.2 428.86 110.06 429.36 ;
      RECT 7.2 430.56 110.06 431.06 ;
      RECT 109.46 430.26 110.06 431.06 ;
      RECT 109.46 432.26 110.06 433.07 ;
      RECT 7.2 432.26 110.06 432.76 ;
      RECT 7.2 433.96 110.06 434.46 ;
      RECT 109.46 433.65 110.06 434.46 ;
      RECT 109.46 435.66 110.06 436.46 ;
      RECT 7.2 435.66 110.06 436.16 ;
      RECT 7.2 437.36 110.06 437.86 ;
      RECT 109.46 437.06 110.06 437.86 ;
      RECT 109.46 439.06 110.06 439.87 ;
      RECT 7.2 439.06 110.06 439.56 ;
      RECT 7.2 440.76 110.06 441.26 ;
      RECT 109.46 440.45 110.06 441.26 ;
      RECT 109.46 442.46 110.06 443.26 ;
      RECT 7.2 442.46 110.06 442.96 ;
      RECT 7.2 444.16 110.06 444.66 ;
      RECT 109.46 443.86 110.06 444.66 ;
      RECT 109.46 445.86 110.06 446.67 ;
      RECT 7.2 445.86 110.06 446.36 ;
      RECT 7.2 447.56 110.06 448.06 ;
      RECT 109.46 447.25 110.06 448.06 ;
      RECT 109.46 449.26 110.06 450.06 ;
      RECT 7.2 449.26 110.06 449.76 ;
      RECT 7.2 450.96 110.06 451.46 ;
      RECT 109.46 450.66 110.06 451.46 ;
      RECT 109.46 452.66 110.06 453.47 ;
      RECT 7.2 452.66 110.06 453.16 ;
      RECT 7.2 454.36 110.06 454.86 ;
      RECT 109.46 454.05 110.06 454.86 ;
      RECT 109.46 456.06 110.06 456.86 ;
      RECT 7.2 456.06 110.06 456.56 ;
      RECT 7.2 457.76 110.06 458.26 ;
      RECT 109.46 457.46 110.06 458.26 ;
      RECT 109.46 459.46 110.06 460.27 ;
      RECT 7.2 459.46 110.06 459.96 ;
      RECT 7.2 461.16 110.06 461.66 ;
      RECT 109.46 460.85 110.06 461.66 ;
      RECT 109.46 462.86 110.06 463.66 ;
      RECT 7.2 462.86 110.06 463.36 ;
      RECT 7.2 464.56 110.06 465.06 ;
      RECT 109.46 464.26 110.06 465.06 ;
      RECT 109.46 466.26 110.06 467.07 ;
      RECT 7.2 466.26 110.06 466.76 ;
      RECT 7.2 467.96 110.06 468.46 ;
      RECT 109.46 467.65 110.06 468.46 ;
      RECT 109.46 469.66 110.06 470.46 ;
      RECT 7.2 469.66 110.06 470.16 ;
      RECT 7.2 471.36 110.06 471.86 ;
      RECT 109.46 471.06 110.06 471.86 ;
      RECT 109.46 473.06 110.06 473.87 ;
      RECT 7.2 473.06 110.06 473.56 ;
      RECT 7.2 474.76 110.06 475.26 ;
      RECT 109.46 474.45 110.06 475.26 ;
      RECT 109.46 476.46 110.06 477.26 ;
      RECT 7.2 476.46 110.06 476.96 ;
      RECT 7.2 478.16 110.06 478.66 ;
      RECT 109.46 477.86 110.06 478.66 ;
      RECT 109.46 479.86 110.06 480.67 ;
      RECT 7.2 479.86 110.06 480.36 ;
      RECT 7.2 481.56 110.06 482.06 ;
      RECT 109.46 481.25 110.06 482.06 ;
      RECT 109.46 483.26 110.06 484.06 ;
      RECT 7.2 483.26 110.06 483.76 ;
      RECT 7.2 484.96 110.06 485.46 ;
      RECT 109.46 484.66 110.06 485.46 ;
      RECT 109.46 486.66 110.06 487.47 ;
      RECT 7.2 486.66 110.06 487.16 ;
      RECT 7.2 488.36 110.06 488.86 ;
      RECT 109.46 488.05 110.06 488.86 ;
      RECT 109.46 490.06 110.06 490.86 ;
      RECT 7.2 490.06 110.06 490.56 ;
      RECT 7.2 491.76 110.06 492.26 ;
      RECT 109.46 491.46 110.06 492.26 ;
      RECT 109.46 493.46 110.06 494.27 ;
      RECT 7.2 493.46 110.06 493.96 ;
      RECT 7.2 495.16 110.06 495.66 ;
      RECT 109.46 494.85 110.06 495.66 ;
      RECT 109.46 496.86 110.06 497.66 ;
      RECT 7.2 496.86 110.06 497.36 ;
      RECT 7.2 498.56 110.06 499.06 ;
      RECT 109.46 498.26 110.06 499.06 ;
      RECT 109.46 500.26 110.06 501.07 ;
      RECT 7.2 500.26 110.06 500.76 ;
      RECT 7.2 501.96 110.06 502.46 ;
      RECT 109.46 501.65 110.06 502.46 ;
      RECT 109.46 503.66 110.06 504.46 ;
      RECT 7.2 503.66 110.06 504.16 ;
      RECT 45.6 508.1 88.1 508.6 ;
      RECT 45.6 506.4 46.1 508.6 ;
      RECT 45.6 506.4 110.06 506.9 ;
      RECT 109.46 505.12 110.06 506.9 ;
      RECT 0 69.16 6.84 69.96 ;
      RECT 0 69.36 88.41 69.76 ;
      RECT 87.83 68.43 88.2 69.76 ;
      RECT 87.83 68.43 109.99 68.63 ;
      RECT 109.39 68.13 109.99 68.63 ;
      RECT 88.41 68.83 88.76 69.16 ;
      RECT 88.41 68.83 109.99 69.03 ;
      RECT 109.36 71.06 109.96 71.56 ;
      RECT 89.86 71.06 109.96 71.46 ;
      RECT 106.16 74.46 109.96 74.86 ;
      RECT 109.36 74.36 109.96 74.86 ;
      RECT 109.36 77.86 109.96 78.36 ;
      RECT 106.16 77.86 109.96 78.26 ;
      RECT 106.16 81.26 109.96 81.66 ;
      RECT 109.36 81.16 109.96 81.66 ;
      RECT 109.36 84.66 109.96 85.16 ;
      RECT 106.16 84.66 109.96 85.06 ;
      RECT 106.16 88.06 109.96 88.46 ;
      RECT 109.36 87.96 109.96 88.46 ;
      RECT 109.36 91.46 109.96 91.96 ;
      RECT 106.16 91.46 109.96 91.86 ;
      RECT 106.16 94.86 109.96 95.26 ;
      RECT 109.36 94.76 109.96 95.26 ;
      RECT 109.36 98.26 109.96 98.76 ;
      RECT 106.16 98.26 109.96 98.66 ;
      RECT 106.16 101.66 109.96 102.06 ;
      RECT 109.36 101.56 109.96 102.06 ;
      RECT 109.36 105.06 109.96 105.56 ;
      RECT 106.16 105.06 109.96 105.46 ;
      RECT 106.16 108.46 109.96 108.86 ;
      RECT 109.36 108.36 109.96 108.86 ;
      RECT 109.36 111.86 109.96 112.36 ;
      RECT 106.16 111.86 109.96 112.26 ;
      RECT 106.16 115.26 109.96 115.66 ;
      RECT 109.36 115.16 109.96 115.66 ;
      RECT 109.36 118.66 109.96 119.16 ;
      RECT 106.16 118.66 109.96 119.06 ;
      RECT 106.16 122.06 109.96 122.46 ;
      RECT 109.36 121.96 109.96 122.46 ;
      RECT 109.36 125.46 109.96 125.96 ;
      RECT 106.16 125.46 109.96 125.86 ;
      RECT 106.16 128.86 109.96 129.26 ;
      RECT 109.36 128.76 109.96 129.26 ;
      RECT 109.36 132.26 109.96 132.76 ;
      RECT 106.16 132.26 109.96 132.66 ;
      RECT 106.16 135.66 109.96 136.06 ;
      RECT 109.36 135.56 109.96 136.06 ;
      RECT 109.36 139.06 109.96 139.56 ;
      RECT 106.16 139.06 109.96 139.46 ;
      RECT 106.16 142.46 109.96 142.86 ;
      RECT 109.36 142.36 109.96 142.86 ;
      RECT 109.36 145.86 109.96 146.36 ;
      RECT 106.16 145.86 109.96 146.26 ;
      RECT 106.16 149.26 109.96 149.66 ;
      RECT 109.36 149.16 109.96 149.66 ;
      RECT 109.36 152.66 109.96 153.16 ;
      RECT 106.16 152.66 109.96 153.06 ;
      RECT 106.16 156.06 109.96 156.46 ;
      RECT 109.36 155.96 109.96 156.46 ;
      RECT 109.36 159.46 109.96 159.96 ;
      RECT 106.16 159.46 109.96 159.86 ;
      RECT 106.16 162.86 109.96 163.26 ;
      RECT 109.36 162.76 109.96 163.26 ;
      RECT 109.36 166.26 109.96 166.76 ;
      RECT 106.16 166.26 109.96 166.66 ;
      RECT 106.16 169.66 109.96 170.06 ;
      RECT 109.36 169.56 109.96 170.06 ;
      RECT 109.36 173.06 109.96 173.56 ;
      RECT 106.16 173.06 109.96 173.46 ;
      RECT 106.16 176.46 109.96 176.86 ;
      RECT 109.36 176.36 109.96 176.86 ;
      RECT 109.36 179.86 109.96 180.36 ;
      RECT 89.86 179.86 109.96 180.26 ;
      RECT 106.16 183.26 109.96 183.66 ;
      RECT 109.36 183.16 109.96 183.66 ;
      RECT 109.36 186.66 109.96 187.16 ;
      RECT 106.16 186.66 109.96 187.06 ;
      RECT 106.16 190.06 109.96 190.46 ;
      RECT 109.36 189.96 109.96 190.46 ;
      RECT 109.36 193.46 109.96 193.96 ;
      RECT 106.16 193.46 109.96 193.86 ;
      RECT 106.16 196.86 109.96 197.26 ;
      RECT 109.36 196.76 109.96 197.26 ;
      RECT 109.36 200.26 109.96 200.76 ;
      RECT 106.16 200.26 109.96 200.66 ;
      RECT 106.16 203.66 109.96 204.06 ;
      RECT 109.36 203.56 109.96 204.06 ;
      RECT 109.36 207.06 109.96 207.56 ;
      RECT 106.16 207.06 109.96 207.46 ;
      RECT 106.16 210.46 109.96 210.86 ;
      RECT 109.36 210.36 109.96 210.86 ;
      RECT 109.36 213.86 109.96 214.36 ;
      RECT 106.16 213.86 109.96 214.26 ;
      RECT 106.16 217.26 109.96 217.66 ;
      RECT 109.36 217.16 109.96 217.66 ;
      RECT 109.36 220.66 109.96 221.16 ;
      RECT 106.16 220.66 109.96 221.06 ;
      RECT 106.16 224.06 109.96 224.46 ;
      RECT 109.36 223.96 109.96 224.46 ;
      RECT 109.36 227.46 109.96 227.96 ;
      RECT 106.16 227.46 109.96 227.86 ;
      RECT 106.16 230.86 109.96 231.26 ;
      RECT 109.36 230.76 109.96 231.26 ;
      RECT 109.36 234.26 109.96 234.76 ;
      RECT 106.16 234.26 109.96 234.66 ;
      RECT 106.16 237.66 109.96 238.06 ;
      RECT 109.36 237.56 109.96 238.06 ;
      RECT 109.36 241.06 109.96 241.56 ;
      RECT 106.16 241.06 109.96 241.46 ;
      RECT 106.16 244.46 109.96 244.86 ;
      RECT 109.36 244.36 109.96 244.86 ;
      RECT 109.36 247.86 109.96 248.36 ;
      RECT 106.16 247.86 109.96 248.26 ;
      RECT 106.16 251.26 109.96 251.66 ;
      RECT 109.36 251.16 109.96 251.66 ;
      RECT 109.36 254.66 109.96 255.16 ;
      RECT 106.16 254.66 109.96 255.06 ;
      RECT 106.16 258.06 109.96 258.46 ;
      RECT 109.36 257.96 109.96 258.46 ;
      RECT 109.36 261.46 109.96 261.96 ;
      RECT 106.16 261.46 109.96 261.86 ;
      RECT 106.16 264.86 109.96 265.26 ;
      RECT 109.36 264.76 109.96 265.26 ;
      RECT 109.36 268.26 109.96 268.76 ;
      RECT 106.16 268.26 109.96 268.66 ;
      RECT 106.16 271.66 109.96 272.06 ;
      RECT 109.36 271.56 109.96 272.06 ;
      RECT 109.36 275.06 109.96 275.56 ;
      RECT 106.16 275.06 109.96 275.46 ;
      RECT 106.16 278.46 109.96 278.86 ;
      RECT 109.36 278.36 109.96 278.86 ;
      RECT 109.36 281.86 109.96 282.36 ;
      RECT 106.16 281.86 109.96 282.26 ;
      RECT 106.16 285.26 109.96 285.66 ;
      RECT 109.36 285.16 109.96 285.66 ;
      RECT 109.36 288.66 109.96 289.16 ;
      RECT 89.86 288.66 109.96 289.06 ;
      RECT 106.16 292.06 109.96 292.46 ;
      RECT 109.36 291.96 109.96 292.46 ;
      RECT 109.36 295.46 109.96 295.96 ;
      RECT 106.16 295.46 109.96 295.86 ;
      RECT 106.16 298.86 109.96 299.26 ;
      RECT 109.36 298.76 109.96 299.26 ;
      RECT 109.36 302.26 109.96 302.76 ;
      RECT 106.16 302.26 109.96 302.66 ;
      RECT 106.16 305.66 109.96 306.06 ;
      RECT 109.36 305.56 109.96 306.06 ;
      RECT 109.36 309.06 109.96 309.56 ;
      RECT 106.16 309.06 109.96 309.46 ;
      RECT 106.16 312.46 109.96 312.86 ;
      RECT 109.36 312.36 109.96 312.86 ;
      RECT 109.36 315.86 109.96 316.36 ;
      RECT 106.16 315.86 109.96 316.26 ;
      RECT 106.16 319.26 109.96 319.66 ;
      RECT 109.36 319.16 109.96 319.66 ;
      RECT 109.36 322.66 109.96 323.16 ;
      RECT 106.16 322.66 109.96 323.06 ;
      RECT 106.16 326.06 109.96 326.46 ;
      RECT 109.36 325.96 109.96 326.46 ;
      RECT 109.36 329.46 109.96 329.96 ;
      RECT 106.16 329.46 109.96 329.86 ;
      RECT 106.16 332.86 109.96 333.26 ;
      RECT 109.36 332.76 109.96 333.26 ;
      RECT 109.36 336.26 109.96 336.76 ;
      RECT 106.16 336.26 109.96 336.66 ;
      RECT 106.16 339.66 109.96 340.06 ;
      RECT 109.36 339.56 109.96 340.06 ;
      RECT 109.36 343.06 109.96 343.56 ;
      RECT 106.16 343.06 109.96 343.46 ;
      RECT 106.16 346.46 109.96 346.86 ;
      RECT 109.36 346.36 109.96 346.86 ;
      RECT 109.36 349.86 109.96 350.36 ;
      RECT 106.16 349.86 109.96 350.26 ;
      RECT 106.16 353.26 109.96 353.66 ;
      RECT 109.36 353.16 109.96 353.66 ;
      RECT 109.36 356.66 109.96 357.16 ;
      RECT 106.16 356.66 109.96 357.06 ;
      RECT 106.16 360.06 109.96 360.46 ;
      RECT 109.36 359.96 109.96 360.46 ;
      RECT 109.36 363.46 109.96 363.96 ;
      RECT 106.16 363.46 109.96 363.86 ;
      RECT 106.16 366.86 109.96 367.26 ;
      RECT 109.36 366.76 109.96 367.26 ;
      RECT 109.36 370.26 109.96 370.76 ;
      RECT 106.16 370.26 109.96 370.66 ;
      RECT 106.16 373.66 109.96 374.06 ;
      RECT 109.36 373.56 109.96 374.06 ;
      RECT 109.36 377.06 109.96 377.56 ;
      RECT 106.16 377.06 109.96 377.46 ;
      RECT 106.16 380.46 109.96 380.86 ;
      RECT 109.36 380.36 109.96 380.86 ;
      RECT 109.36 383.86 109.96 384.36 ;
      RECT 106.16 383.86 109.96 384.26 ;
      RECT 106.16 387.26 109.96 387.66 ;
      RECT 109.36 387.16 109.96 387.66 ;
      RECT 109.36 390.66 109.96 391.16 ;
      RECT 106.16 390.66 109.96 391.06 ;
      RECT 106.16 394.06 109.96 394.46 ;
      RECT 109.36 393.96 109.96 394.46 ;
      RECT 109.36 397.46 109.96 397.96 ;
      RECT 89.86 397.46 109.96 397.86 ;
      RECT 106.16 400.86 109.96 401.26 ;
      RECT 109.36 400.76 109.96 401.26 ;
      RECT 109.36 404.26 109.96 404.76 ;
      RECT 106.16 404.26 109.96 404.66 ;
      RECT 106.16 407.66 109.96 408.06 ;
      RECT 109.36 407.56 109.96 408.06 ;
      RECT 109.36 411.06 109.96 411.56 ;
      RECT 106.16 411.06 109.96 411.46 ;
      RECT 106.16 414.46 109.96 414.86 ;
      RECT 109.36 414.36 109.96 414.86 ;
      RECT 109.36 417.86 109.96 418.36 ;
      RECT 106.16 417.86 109.96 418.26 ;
      RECT 106.16 421.26 109.96 421.66 ;
      RECT 109.36 421.16 109.96 421.66 ;
      RECT 109.36 424.66 109.96 425.16 ;
      RECT 106.16 424.66 109.96 425.06 ;
      RECT 106.16 428.06 109.96 428.46 ;
      RECT 109.36 427.96 109.96 428.46 ;
      RECT 109.36 431.46 109.96 431.96 ;
      RECT 106.16 431.46 109.96 431.86 ;
      RECT 106.16 434.86 109.96 435.26 ;
      RECT 109.36 434.76 109.96 435.26 ;
      RECT 109.36 438.26 109.96 438.76 ;
      RECT 106.16 438.26 109.96 438.66 ;
      RECT 106.16 441.66 109.96 442.06 ;
      RECT 109.36 441.56 109.96 442.06 ;
      RECT 109.36 445.06 109.96 445.56 ;
      RECT 106.16 445.06 109.96 445.46 ;
      RECT 106.16 448.46 109.96 448.86 ;
      RECT 109.36 448.36 109.96 448.86 ;
      RECT 109.36 451.86 109.96 452.36 ;
      RECT 106.16 451.86 109.96 452.26 ;
      RECT 106.16 455.26 109.96 455.66 ;
      RECT 109.36 455.16 109.96 455.66 ;
      RECT 109.36 458.66 109.96 459.16 ;
      RECT 106.16 458.66 109.96 459.06 ;
      RECT 106.16 462.06 109.96 462.46 ;
      RECT 109.36 461.96 109.96 462.46 ;
      RECT 109.36 465.46 109.96 465.96 ;
      RECT 106.16 465.46 109.96 465.86 ;
      RECT 106.16 468.86 109.96 469.26 ;
      RECT 109.36 468.76 109.96 469.26 ;
      RECT 109.36 472.26 109.96 472.76 ;
      RECT 106.16 472.26 109.96 472.66 ;
      RECT 106.16 475.66 109.96 476.06 ;
      RECT 109.36 475.56 109.96 476.06 ;
      RECT 109.36 479.06 109.96 479.56 ;
      RECT 106.16 479.06 109.96 479.46 ;
      RECT 106.16 482.46 109.96 482.86 ;
      RECT 109.36 482.36 109.96 482.86 ;
      RECT 109.36 485.86 109.96 486.36 ;
      RECT 106.16 485.86 109.96 486.26 ;
      RECT 106.16 489.26 109.96 489.66 ;
      RECT 109.36 489.16 109.96 489.66 ;
      RECT 109.36 492.66 109.96 493.16 ;
      RECT 106.16 492.66 109.96 493.06 ;
      RECT 106.16 496.06 109.96 496.46 ;
      RECT 109.36 495.96 109.96 496.46 ;
      RECT 109.36 499.46 109.96 499.96 ;
      RECT 106.16 499.46 109.96 499.86 ;
      RECT 106.16 502.86 109.96 503.26 ;
      RECT 109.36 502.76 109.96 503.26 ;
      RECT 107.63 66.03 108.13 66.43 ;
      RECT 107.83 54.14 108.13 66.43 ;
      RECT 107.41 54.14 108.13 54.44 ;
      RECT 107.41 44.24 107.71 54.44 ;
      RECT 107.41 16.13 107.61 54.44 ;
      RECT 106.86 65.53 107.34 66.43 ;
      RECT 106.86 65.53 107.61 65.83 ;
      RECT 107.41 61.91 107.61 65.83 ;
      RECT 105.31 39.44 106.31 66.63 ;
      RECT 105.61 6.24 106.01 66.63 ;
      RECT 104.83 6.24 106.79 32.15 ;
      RECT 104.92 34.93 105.12 38.18 ;
      RECT 104.41 34.93 105.12 35.13 ;
      RECT 104.41 12.32 104.61 35.13 ;
      RECT 104.24 66.04 104.89 66.43 ;
      RECT 104.59 61.1 104.89 66.43 ;
      RECT 103.92 61.1 104.89 61.4 ;
      RECT 103.92 44.24 104.22 61.4 ;
      RECT 104.01 16.13 104.21 61.4 ;
      RECT 103.46 65.53 103.94 66.43 ;
      RECT 103.46 65.53 104.21 65.83 ;
      RECT 104.01 61.91 104.21 65.83 ;
      RECT 101.91 39.44 102.91 66.63 ;
      RECT 102.21 6.24 102.61 66.63 ;
      RECT 101.43 6.24 103.39 32.15 ;
      RECT 100.83 66.03 101.33 66.43 ;
      RECT 101.03 54.14 101.33 66.43 ;
      RECT 100.61 54.14 101.33 54.44 ;
      RECT 100.61 44.24 100.91 54.44 ;
      RECT 100.61 16.13 100.81 54.44 ;
      RECT 100.06 65.53 100.54 66.43 ;
      RECT 100.06 65.53 100.81 65.83 ;
      RECT 100.61 61.91 100.81 65.83 ;
      RECT 98.51 39.44 99.51 66.63 ;
      RECT 98.81 6.24 99.21 66.63 ;
      RECT 98.01 6.24 99.99 32.15 ;
      RECT 97.43 66.03 98.09 66.43 ;
      RECT 97.79 61.1 98.09 66.43 ;
      RECT 97.12 61.1 98.09 61.4 ;
      RECT 97.12 44.24 97.42 61.4 ;
      RECT 97.21 16.13 97.41 61.4 ;
      RECT 96.66 65.53 97.14 66.43 ;
      RECT 96.66 65.53 97.41 65.83 ;
      RECT 97.21 61.91 97.41 65.83 ;
      RECT 95.41 6.24 95.81 66.63 ;
      RECT 95.11 6.24 95.81 54.64 ;
      RECT 95.11 39.44 96.11 54.42 ;
      RECT 95.11 6.24 96.61 32.15 ;
      RECT 94.63 6.24 96.61 15.28 ;
      RECT 94.04 65.63 94.51 66.33 ;
      RECT 93.73 65.63 94.51 65.83 ;
      RECT 93.81 61.91 94.01 65.83 ;
      RECT 93.26 66.03 93.74 66.33 ;
      RECT 93.26 60.97 93.46 66.33 ;
      RECT 93.26 60.97 94.01 61.17 ;
      RECT 93.81 16.13 94.01 61.17 ;
      RECT 92.01 6.24 92.41 66.63 ;
      RECT 91.71 40.16 92.71 65.02 ;
      RECT 91.71 6.24 92.71 31.95 ;
      RECT 91.23 6.24 93.19 15.28 ;
      RECT 91.32 35.33 91.52 38.18 ;
      RECT 90.81 35.33 91.52 35.53 ;
      RECT 90.81 12.32 91.01 35.53 ;
      RECT 90.64 65.63 91.11 66.33 ;
      RECT 90.41 65.63 91.11 65.83 ;
      RECT 90.41 61.91 90.61 65.83 ;
      RECT 89.86 66.03 90.34 66.33 ;
      RECT 89.86 54.04 90.06 66.33 ;
      RECT 89.86 54.04 90.61 54.24 ;
      RECT 90.41 16.13 90.61 54.24 ;
      RECT 88.61 6.24 89.01 66.63 ;
      RECT 88.61 6.24 89.31 54.64 ;
      RECT 88.61 6.24 89.79 15.28 ;
      RECT 0 72.56 6.84 73.36 ;
      RECT 0 72.76 88.61 73.16 ;
      RECT 0 79.36 6.84 80.16 ;
      RECT 0 79.56 88.61 79.96 ;
      RECT 0 86.16 6.84 86.96 ;
      RECT 0 86.36 88.61 86.76 ;
      RECT 0 92.96 6.84 93.76 ;
      RECT 0 93.16 88.61 93.56 ;
      RECT 0 99.76 6.84 100.56 ;
      RECT 0 99.96 88.61 100.36 ;
      RECT 0 106.56 6.84 107.36 ;
      RECT 0 106.76 88.61 107.16 ;
      RECT 0 113.36 6.84 114.16 ;
      RECT 0 113.56 88.61 113.96 ;
      RECT 0 120.16 6.84 120.96 ;
      RECT 0 120.36 88.61 120.76 ;
      RECT 0 126.96 6.84 127.76 ;
      RECT 0 127.16 88.61 127.56 ;
      RECT 0 133.76 6.84 134.56 ;
      RECT 0 133.96 88.61 134.36 ;
      RECT 0 140.56 6.84 141.36 ;
      RECT 0 140.76 88.61 141.16 ;
      RECT 0 147.36 6.84 148.16 ;
      RECT 0 147.56 88.61 147.96 ;
      RECT 0 154.16 6.84 154.96 ;
      RECT 0 154.36 88.61 154.76 ;
      RECT 0 160.96 6.84 161.76 ;
      RECT 0 161.16 88.61 161.56 ;
      RECT 0 167.76 6.84 168.56 ;
      RECT 0 167.96 88.61 168.36 ;
      RECT 0 174.56 6.84 175.36 ;
      RECT 0 174.76 88.61 175.16 ;
      RECT 0 181.36 6.84 182.16 ;
      RECT 0 181.56 88.61 181.96 ;
      RECT 0 188.16 6.84 188.96 ;
      RECT 0 188.36 88.61 188.76 ;
      RECT 0 194.96 6.84 195.76 ;
      RECT 0 195.16 88.61 195.56 ;
      RECT 0 201.76 6.84 202.56 ;
      RECT 0 201.96 88.61 202.36 ;
      RECT 0 208.56 6.84 209.36 ;
      RECT 0 208.76 88.61 209.16 ;
      RECT 0 215.36 6.84 216.16 ;
      RECT 0 215.56 88.61 215.96 ;
      RECT 0 222.16 6.84 222.96 ;
      RECT 0 222.36 88.61 222.76 ;
      RECT 0 228.96 6.84 229.76 ;
      RECT 0 229.16 88.61 229.56 ;
      RECT 0 235.76 6.84 236.56 ;
      RECT 0 235.96 88.61 236.36 ;
      RECT 0 242.56 6.84 243.36 ;
      RECT 0 242.76 88.61 243.16 ;
      RECT 0 249.36 6.84 250.16 ;
      RECT 0 249.56 88.61 249.96 ;
      RECT 0 256.16 6.84 256.96 ;
      RECT 0 256.36 88.61 256.76 ;
      RECT 0 262.96 6.84 263.76 ;
      RECT 0 263.16 88.61 263.56 ;
      RECT 0 269.76 6.84 270.56 ;
      RECT 0 269.96 88.61 270.36 ;
      RECT 0 276.56 6.84 277.36 ;
      RECT 0 276.76 88.61 277.16 ;
      RECT 0 283.36 6.84 284.16 ;
      RECT 0 283.56 88.61 283.96 ;
      RECT 0 290.16 6.84 290.96 ;
      RECT 0 290.36 88.61 290.76 ;
      RECT 0 296.96 6.84 297.76 ;
      RECT 0 297.16 88.61 297.56 ;
      RECT 0 303.76 6.84 304.56 ;
      RECT 0 303.96 88.61 304.36 ;
      RECT 0 310.56 6.84 311.36 ;
      RECT 0 310.76 88.61 311.16 ;
      RECT 0 317.36 6.84 318.16 ;
      RECT 0 317.56 88.61 317.96 ;
      RECT 0 324.16 6.84 324.96 ;
      RECT 0 324.36 88.61 324.76 ;
      RECT 0 330.96 6.84 331.76 ;
      RECT 0 331.16 88.61 331.56 ;
      RECT 0 337.76 6.84 338.56 ;
      RECT 0 337.96 88.61 338.36 ;
      RECT 0 344.56 6.84 345.36 ;
      RECT 0 344.76 88.61 345.16 ;
      RECT 0 351.36 6.84 352.16 ;
      RECT 0 351.56 88.61 351.96 ;
      RECT 0 358.16 6.84 358.96 ;
      RECT 0 358.36 88.61 358.76 ;
      RECT 0 364.96 6.84 365.76 ;
      RECT 0 365.16 88.61 365.56 ;
      RECT 0 371.76 6.84 372.56 ;
      RECT 0 371.96 88.61 372.36 ;
      RECT 0 378.56 6.84 379.36 ;
      RECT 0 378.76 88.61 379.16 ;
      RECT 0 385.36 6.84 386.16 ;
      RECT 0 385.56 88.61 385.96 ;
      RECT 0 392.16 6.84 392.96 ;
      RECT 0 392.36 88.61 392.76 ;
      RECT 0 398.96 6.84 399.76 ;
      RECT 0 399.16 88.61 399.56 ;
      RECT 0 405.76 6.84 406.56 ;
      RECT 0 405.96 88.61 406.36 ;
      RECT 0 412.56 6.84 413.36 ;
      RECT 0 412.76 88.61 413.16 ;
      RECT 0 419.36 6.84 420.16 ;
      RECT 0 419.56 88.61 419.96 ;
      RECT 0 426.16 6.84 426.96 ;
      RECT 0 426.36 88.61 426.76 ;
      RECT 0 432.96 6.84 433.76 ;
      RECT 0 433.16 88.61 433.56 ;
      RECT 0 439.76 6.84 440.56 ;
      RECT 0 439.96 88.61 440.36 ;
      RECT 0 446.56 6.84 447.36 ;
      RECT 0 446.76 88.61 447.16 ;
      RECT 0 453.36 6.84 454.16 ;
      RECT 0 453.56 88.61 453.96 ;
      RECT 0 460.16 6.84 460.96 ;
      RECT 0 460.36 88.61 460.76 ;
      RECT 0 466.96 6.84 467.76 ;
      RECT 0 467.16 88.61 467.56 ;
      RECT 0 473.76 6.84 474.56 ;
      RECT 0 473.96 88.61 474.36 ;
      RECT 0 480.56 6.84 481.36 ;
      RECT 0 480.76 88.61 481.16 ;
      RECT 0 487.36 6.84 488.16 ;
      RECT 0 487.56 88.61 487.96 ;
      RECT 0 494.16 6.84 494.96 ;
      RECT 0 494.36 88.61 494.76 ;
      RECT 0 500.96 6.84 501.76 ;
      RECT 0 501.16 88.61 501.56 ;
      RECT 0 75.96 6.84 76.76 ;
      RECT 0 76.16 88.41 76.56 ;
      RECT 0 82.76 6.84 83.56 ;
      RECT 0 82.96 88.41 83.36 ;
      RECT 0 89.56 6.84 90.36 ;
      RECT 0 89.76 88.41 90.16 ;
      RECT 0 96.36 6.84 97.16 ;
      RECT 0 96.56 88.41 96.96 ;
      RECT 0 103.16 6.84 103.96 ;
      RECT 0 103.36 88.41 103.76 ;
      RECT 0 109.96 6.84 110.76 ;
      RECT 0 110.16 88.41 110.56 ;
      RECT 0 116.76 6.84 117.56 ;
      RECT 0 116.96 88.41 117.36 ;
      RECT 0 123.56 6.84 124.36 ;
      RECT 0 123.76 88.41 124.16 ;
      RECT 0 130.36 6.84 131.16 ;
      RECT 0 130.56 88.41 130.96 ;
      RECT 0 137.16 6.84 137.96 ;
      RECT 0 137.36 88.41 137.76 ;
      RECT 0 143.96 6.84 144.76 ;
      RECT 0 144.16 88.41 144.56 ;
      RECT 0 150.76 6.84 151.56 ;
      RECT 0 150.96 88.41 151.36 ;
      RECT 0 157.56 6.84 158.36 ;
      RECT 0 157.76 88.41 158.16 ;
      RECT 0 164.36 6.84 165.16 ;
      RECT 0 164.56 88.41 164.96 ;
      RECT 0 171.16 6.84 171.96 ;
      RECT 0 171.36 88.41 171.76 ;
      RECT 0 177.96 6.84 178.76 ;
      RECT 0 178.16 88.41 178.56 ;
      RECT 0 184.76 6.84 185.56 ;
      RECT 0 184.96 88.41 185.36 ;
      RECT 0 191.56 6.84 192.36 ;
      RECT 0 191.76 88.41 192.16 ;
      RECT 0 198.36 6.84 199.16 ;
      RECT 0 198.56 88.41 198.96 ;
      RECT 0 205.16 6.84 205.96 ;
      RECT 0 205.36 88.41 205.76 ;
      RECT 0 211.96 6.84 212.76 ;
      RECT 0 212.16 88.41 212.56 ;
      RECT 0 218.76 6.84 219.56 ;
      RECT 0 218.96 88.41 219.36 ;
      RECT 0 225.56 6.84 226.36 ;
      RECT 0 225.76 88.41 226.16 ;
      RECT 0 232.36 6.84 233.16 ;
      RECT 0 232.56 88.41 232.96 ;
      RECT 0 239.16 6.84 239.96 ;
      RECT 0 239.36 88.41 239.76 ;
      RECT 0 245.96 6.84 246.76 ;
      RECT 0 246.16 88.41 246.56 ;
      RECT 0 252.76 6.84 253.56 ;
      RECT 0 252.96 88.41 253.36 ;
      RECT 0 259.56 6.84 260.36 ;
      RECT 0 259.76 88.41 260.16 ;
      RECT 0 266.36 6.84 267.16 ;
      RECT 0 266.56 88.41 266.96 ;
      RECT 0 273.16 6.84 273.96 ;
      RECT 0 273.36 88.41 273.76 ;
      RECT 0 279.96 6.84 280.76 ;
      RECT 0 280.16 88.41 280.56 ;
      RECT 0 286.76 6.84 287.56 ;
      RECT 0 286.96 88.41 287.36 ;
      RECT 0 293.56 6.84 294.36 ;
      RECT 0 293.76 88.41 294.16 ;
      RECT 0 300.36 6.84 301.16 ;
      RECT 0 300.56 88.41 300.96 ;
      RECT 0 307.16 6.84 307.96 ;
      RECT 0 307.36 88.41 307.76 ;
      RECT 0 313.96 6.84 314.76 ;
      RECT 0 314.16 88.41 314.56 ;
      RECT 0 320.76 6.84 321.56 ;
      RECT 0 320.96 88.41 321.36 ;
      RECT 0 327.56 6.84 328.36 ;
      RECT 0 327.76 88.41 328.16 ;
      RECT 0 334.36 6.84 335.16 ;
      RECT 0 334.56 88.41 334.96 ;
      RECT 0 341.16 6.84 341.96 ;
      RECT 0 341.36 88.41 341.76 ;
      RECT 0 347.96 6.84 348.76 ;
      RECT 0 348.16 88.41 348.56 ;
      RECT 0 354.76 6.84 355.56 ;
      RECT 0 354.96 88.41 355.36 ;
      RECT 0 361.56 6.84 362.36 ;
      RECT 0 361.76 88.41 362.16 ;
      RECT 0 368.36 6.84 369.16 ;
      RECT 0 368.56 88.41 368.96 ;
      RECT 0 375.16 6.84 375.96 ;
      RECT 0 375.36 88.41 375.76 ;
      RECT 0 381.96 6.84 382.76 ;
      RECT 0 382.16 88.41 382.56 ;
      RECT 0 388.76 6.84 389.56 ;
      RECT 0 388.96 88.41 389.36 ;
      RECT 0 395.56 6.84 396.36 ;
      RECT 0 395.76 88.41 396.16 ;
      RECT 0 402.36 6.84 403.16 ;
      RECT 0 402.56 88.41 402.96 ;
      RECT 0 409.16 6.84 409.96 ;
      RECT 0 409.36 88.41 409.76 ;
      RECT 0 415.96 6.84 416.76 ;
      RECT 0 416.16 88.41 416.56 ;
      RECT 0 422.76 6.84 423.56 ;
      RECT 0 422.96 88.41 423.36 ;
      RECT 0 429.56 6.84 430.36 ;
      RECT 0 429.76 88.41 430.16 ;
      RECT 0 436.36 6.84 437.16 ;
      RECT 0 436.56 88.41 436.96 ;
      RECT 0 443.16 6.84 443.96 ;
      RECT 0 443.36 88.41 443.76 ;
      RECT 0 449.96 6.84 450.76 ;
      RECT 0 450.16 88.41 450.56 ;
      RECT 0 456.76 6.84 457.56 ;
      RECT 0 456.96 88.41 457.36 ;
      RECT 0 463.56 6.84 464.36 ;
      RECT 0 463.76 88.41 464.16 ;
      RECT 0 470.36 6.84 471.16 ;
      RECT 0 470.56 88.41 470.96 ;
      RECT 0 477.16 6.84 477.96 ;
      RECT 0 477.36 88.41 477.76 ;
      RECT 0 483.96 6.84 484.76 ;
      RECT 0 484.16 88.41 484.56 ;
      RECT 0 490.76 6.84 491.56 ;
      RECT 0 490.96 88.41 491.36 ;
      RECT 0 497.56 6.84 498.36 ;
      RECT 0 497.76 88.41 498.16 ;
      RECT 0 504.36 6.84 505.16 ;
      RECT 0 504.56 88.41 504.96 ;
      RECT 83.01 509 85.01 510.94 ;
      RECT 78.21 509 80.21 510.94 ;
      RECT 73.41 509 75.41 510.94 ;
      RECT 68.61 509 70.61 510.94 ;
      RECT 63.81 509 65.81 510.94 ;
      RECT 59.01 509 61.01 510.94 ;
      RECT 54.21 509 56.21 510.94 ;
      RECT 49.41 509 51.41 510.94 ;
      RECT 43.41 509 45.41 510.94 ;
      RECT 38.61 509 40.61 510.94 ;
      RECT 33.81 509 35.81 510.94 ;
      RECT 29.01 509 31.01 510.94 ;
      RECT 24.21 509 26.21 510.94 ;
      RECT 19.41 509 21.41 510.94 ;
      RECT 14.61 509 16.61 510.94 ;
      RECT 9.81 509 11.81 510.94 ;
      RECT 0 509 6.84 509.8 ;
      RECT 0 509 88.2 509.4 ;
      RECT 3.12 70.86 6.84 71.66 ;
      RECT 3.12 71.06 88.1 71.46 ;
      RECT 3.12 74.26 6.84 75.06 ;
      RECT 3.12 74.46 88.1 74.86 ;
      RECT 3.12 77.66 6.84 78.46 ;
      RECT 3.12 77.86 88.1 78.26 ;
      RECT 3.12 81.06 6.84 81.86 ;
      RECT 3.12 81.26 88.1 81.66 ;
      RECT 3.12 84.46 6.84 85.26 ;
      RECT 3.12 84.66 88.1 85.06 ;
      RECT 3.12 87.86 6.84 88.66 ;
      RECT 3.12 88.06 88.1 88.46 ;
      RECT 3.12 91.26 6.84 92.06 ;
      RECT 3.12 91.46 88.1 91.86 ;
      RECT 3.12 94.66 6.84 95.46 ;
      RECT 3.12 94.86 88.1 95.26 ;
      RECT 3.12 98.06 6.84 98.86 ;
      RECT 3.12 98.26 88.1 98.66 ;
      RECT 3.12 101.46 6.84 102.26 ;
      RECT 3.12 101.66 88.1 102.06 ;
      RECT 3.12 104.86 6.84 105.66 ;
      RECT 3.12 105.06 88.1 105.46 ;
      RECT 3.12 108.26 6.84 109.06 ;
      RECT 3.12 108.46 88.1 108.86 ;
      RECT 3.12 111.66 6.84 112.46 ;
      RECT 3.12 111.86 88.1 112.26 ;
      RECT 3.12 115.06 6.84 115.86 ;
      RECT 3.12 115.26 88.1 115.66 ;
      RECT 3.12 118.46 6.84 119.26 ;
      RECT 3.12 118.66 88.1 119.06 ;
      RECT 3.12 121.86 6.84 122.66 ;
      RECT 3.12 122.06 88.1 122.46 ;
      RECT 3.12 125.26 6.84 126.06 ;
      RECT 3.12 125.46 88.1 125.86 ;
      RECT 3.12 128.66 6.84 129.46 ;
      RECT 3.12 128.86 88.1 129.26 ;
      RECT 3.12 132.06 6.84 132.86 ;
      RECT 3.12 132.26 88.1 132.66 ;
      RECT 3.12 135.46 6.84 136.26 ;
      RECT 3.12 135.66 88.1 136.06 ;
      RECT 3.12 138.86 6.84 139.66 ;
      RECT 3.12 139.06 88.1 139.46 ;
      RECT 3.12 142.26 6.84 143.06 ;
      RECT 3.12 142.46 88.1 142.86 ;
      RECT 3.12 145.66 6.84 146.46 ;
      RECT 3.12 145.86 88.1 146.26 ;
      RECT 3.12 149.06 6.84 149.86 ;
      RECT 3.12 149.26 88.1 149.66 ;
      RECT 3.12 152.46 6.84 153.26 ;
      RECT 3.12 152.66 88.1 153.06 ;
      RECT 3.12 155.86 6.84 156.66 ;
      RECT 3.12 156.06 88.1 156.46 ;
      RECT 3.12 159.26 6.84 160.06 ;
      RECT 3.12 159.46 88.1 159.86 ;
      RECT 3.12 162.66 6.84 163.46 ;
      RECT 3.12 162.86 88.1 163.26 ;
      RECT 3.12 166.06 6.84 166.86 ;
      RECT 3.12 166.26 88.1 166.66 ;
      RECT 3.12 169.46 6.84 170.26 ;
      RECT 3.12 169.66 88.1 170.06 ;
      RECT 3.12 172.86 6.84 173.66 ;
      RECT 3.12 173.06 88.1 173.46 ;
      RECT 3.12 176.26 6.84 177.06 ;
      RECT 3.12 176.46 88.1 176.86 ;
      RECT 3.12 179.66 6.84 180.46 ;
      RECT 3.12 179.86 88.1 180.26 ;
      RECT 3.12 183.06 6.84 183.86 ;
      RECT 3.12 183.26 88.1 183.66 ;
      RECT 3.12 186.46 6.84 187.26 ;
      RECT 3.12 186.66 88.1 187.06 ;
      RECT 3.12 189.86 6.84 190.66 ;
      RECT 3.12 190.06 88.1 190.46 ;
      RECT 3.12 193.26 6.84 194.06 ;
      RECT 3.12 193.46 88.1 193.86 ;
      RECT 3.12 196.66 6.84 197.46 ;
      RECT 3.12 196.86 88.1 197.26 ;
      RECT 3.12 200.06 6.84 200.86 ;
      RECT 3.12 200.26 88.1 200.66 ;
      RECT 3.12 203.46 6.84 204.26 ;
      RECT 3.12 203.66 88.1 204.06 ;
      RECT 3.12 206.86 6.84 207.66 ;
      RECT 3.12 207.06 88.1 207.46 ;
      RECT 3.12 210.26 6.84 211.06 ;
      RECT 3.12 210.46 88.1 210.86 ;
      RECT 3.12 213.66 6.84 214.46 ;
      RECT 3.12 213.86 88.1 214.26 ;
      RECT 3.12 217.06 6.84 217.86 ;
      RECT 3.12 217.26 88.1 217.66 ;
      RECT 3.12 220.46 6.84 221.26 ;
      RECT 3.12 220.66 88.1 221.06 ;
      RECT 3.12 223.86 6.84 224.66 ;
      RECT 3.12 224.06 88.1 224.46 ;
      RECT 3.12 227.26 6.84 228.06 ;
      RECT 3.12 227.46 88.1 227.86 ;
      RECT 3.12 230.66 6.84 231.46 ;
      RECT 3.12 230.86 88.1 231.26 ;
      RECT 3.12 234.06 6.84 234.86 ;
      RECT 3.12 234.26 88.1 234.66 ;
      RECT 3.12 237.46 6.84 238.26 ;
      RECT 3.12 237.66 88.1 238.06 ;
      RECT 3.12 240.86 6.84 241.66 ;
      RECT 3.12 241.06 88.1 241.46 ;
      RECT 3.12 244.26 6.84 245.06 ;
      RECT 3.12 244.46 88.1 244.86 ;
      RECT 3.12 247.66 6.84 248.46 ;
      RECT 3.12 247.86 88.1 248.26 ;
      RECT 3.12 251.06 6.84 251.86 ;
      RECT 3.12 251.26 88.1 251.66 ;
      RECT 3.12 254.46 6.84 255.26 ;
      RECT 3.12 254.66 88.1 255.06 ;
      RECT 3.12 257.86 6.84 258.66 ;
      RECT 3.12 258.06 88.1 258.46 ;
      RECT 3.12 261.26 6.84 262.06 ;
      RECT 3.12 261.46 88.1 261.86 ;
      RECT 3.12 264.66 6.84 265.46 ;
      RECT 3.12 264.86 88.1 265.26 ;
      RECT 3.12 268.06 6.84 268.86 ;
      RECT 3.12 268.26 88.1 268.66 ;
      RECT 3.12 271.46 6.84 272.26 ;
      RECT 3.12 271.66 88.1 272.06 ;
      RECT 3.12 274.86 6.84 275.66 ;
      RECT 3.12 275.06 88.1 275.46 ;
      RECT 3.12 278.26 6.84 279.06 ;
      RECT 3.12 278.46 88.1 278.86 ;
      RECT 3.12 281.66 6.84 282.46 ;
      RECT 3.12 281.86 88.1 282.26 ;
      RECT 3.12 285.06 6.84 285.86 ;
      RECT 3.12 285.26 88.1 285.66 ;
      RECT 3.12 288.46 6.84 289.26 ;
      RECT 3.12 288.66 88.1 289.06 ;
      RECT 3.12 291.86 6.84 292.66 ;
      RECT 3.12 292.06 88.1 292.46 ;
      RECT 3.12 295.26 6.84 296.06 ;
      RECT 3.12 295.46 88.1 295.86 ;
      RECT 3.12 298.66 6.84 299.46 ;
      RECT 3.12 298.86 88.1 299.26 ;
      RECT 3.12 302.06 6.84 302.86 ;
      RECT 3.12 302.26 88.1 302.66 ;
      RECT 3.12 305.46 6.84 306.26 ;
      RECT 3.12 305.66 88.1 306.06 ;
      RECT 3.12 308.86 6.84 309.66 ;
      RECT 3.12 309.06 88.1 309.46 ;
      RECT 3.12 312.26 6.84 313.06 ;
      RECT 3.12 312.46 88.1 312.86 ;
      RECT 3.12 315.66 6.84 316.46 ;
      RECT 3.12 315.86 88.1 316.26 ;
      RECT 3.12 319.06 6.84 319.86 ;
      RECT 3.12 319.26 88.1 319.66 ;
      RECT 3.12 322.46 6.84 323.26 ;
      RECT 3.12 322.66 88.1 323.06 ;
      RECT 3.12 325.86 6.84 326.66 ;
      RECT 3.12 326.06 88.1 326.46 ;
      RECT 3.12 329.26 6.84 330.06 ;
      RECT 3.12 329.46 88.1 329.86 ;
      RECT 3.12 332.66 6.84 333.46 ;
      RECT 3.12 332.86 88.1 333.26 ;
      RECT 3.12 336.06 6.84 336.86 ;
      RECT 3.12 336.26 88.1 336.66 ;
      RECT 3.12 339.46 6.84 340.26 ;
      RECT 3.12 339.66 88.1 340.06 ;
      RECT 3.12 342.86 6.84 343.66 ;
      RECT 3.12 343.06 88.1 343.46 ;
      RECT 3.12 346.26 6.84 347.06 ;
      RECT 3.12 346.46 88.1 346.86 ;
      RECT 3.12 349.66 6.84 350.46 ;
      RECT 3.12 349.86 88.1 350.26 ;
      RECT 3.12 353.06 6.84 353.86 ;
      RECT 3.12 353.26 88.1 353.66 ;
      RECT 3.12 356.46 6.84 357.26 ;
      RECT 3.12 356.66 88.1 357.06 ;
      RECT 3.12 359.86 6.84 360.66 ;
      RECT 3.12 360.06 88.1 360.46 ;
      RECT 3.12 363.26 6.84 364.06 ;
      RECT 3.12 363.46 88.1 363.86 ;
      RECT 3.12 366.66 6.84 367.46 ;
      RECT 3.12 366.86 88.1 367.26 ;
      RECT 3.12 370.06 6.84 370.86 ;
      RECT 3.12 370.26 88.1 370.66 ;
      RECT 3.12 373.46 6.84 374.26 ;
      RECT 3.12 373.66 88.1 374.06 ;
      RECT 3.12 376.86 6.84 377.66 ;
      RECT 3.12 377.06 88.1 377.46 ;
      RECT 3.12 380.26 6.84 381.06 ;
      RECT 3.12 380.46 88.1 380.86 ;
      RECT 3.12 383.66 6.84 384.46 ;
      RECT 3.12 383.86 88.1 384.26 ;
      RECT 3.12 387.06 6.84 387.86 ;
      RECT 3.12 387.26 88.1 387.66 ;
      RECT 3.12 390.46 6.84 391.26 ;
      RECT 3.12 390.66 88.1 391.06 ;
      RECT 3.12 393.86 6.84 394.66 ;
      RECT 3.12 394.06 88.1 394.46 ;
      RECT 3.12 397.26 6.84 398.06 ;
      RECT 3.12 397.46 88.1 397.86 ;
      RECT 3.12 400.66 6.84 401.46 ;
      RECT 3.12 400.86 88.1 401.26 ;
      RECT 3.12 404.06 6.84 404.86 ;
      RECT 3.12 404.26 88.1 404.66 ;
      RECT 3.12 407.46 6.84 408.26 ;
      RECT 3.12 407.66 88.1 408.06 ;
      RECT 3.12 410.86 6.84 411.66 ;
      RECT 3.12 411.06 88.1 411.46 ;
      RECT 3.12 414.26 6.84 415.06 ;
      RECT 3.12 414.46 88.1 414.86 ;
      RECT 3.12 417.66 6.84 418.46 ;
      RECT 3.12 417.86 88.1 418.26 ;
      RECT 3.12 421.06 6.84 421.86 ;
      RECT 3.12 421.26 88.1 421.66 ;
      RECT 3.12 424.46 6.84 425.26 ;
      RECT 3.12 424.66 88.1 425.06 ;
      RECT 3.12 427.86 6.84 428.66 ;
      RECT 3.12 428.06 88.1 428.46 ;
      RECT 3.12 431.26 6.84 432.06 ;
      RECT 3.12 431.46 88.1 431.86 ;
      RECT 3.12 434.66 6.84 435.46 ;
      RECT 3.12 434.86 88.1 435.26 ;
      RECT 3.12 438.06 6.84 438.86 ;
      RECT 3.12 438.26 88.1 438.66 ;
      RECT 3.12 441.46 6.84 442.26 ;
      RECT 3.12 441.66 88.1 442.06 ;
      RECT 3.12 444.86 6.84 445.66 ;
      RECT 3.12 445.06 88.1 445.46 ;
      RECT 3.12 448.26 6.84 449.06 ;
      RECT 3.12 448.46 88.1 448.86 ;
      RECT 3.12 451.66 6.84 452.46 ;
      RECT 3.12 451.86 88.1 452.26 ;
      RECT 3.12 455.06 6.84 455.86 ;
      RECT 3.12 455.26 88.1 455.66 ;
      RECT 3.12 458.46 6.84 459.26 ;
      RECT 3.12 458.66 88.1 459.06 ;
      RECT 3.12 461.86 6.84 462.66 ;
      RECT 3.12 462.06 88.1 462.46 ;
      RECT 3.12 465.26 6.84 466.06 ;
      RECT 3.12 465.46 88.1 465.86 ;
      RECT 3.12 468.66 6.84 469.46 ;
      RECT 3.12 468.86 88.1 469.26 ;
      RECT 3.12 472.06 6.84 472.86 ;
      RECT 3.12 472.26 88.1 472.66 ;
      RECT 3.12 475.46 6.84 476.26 ;
      RECT 3.12 475.66 88.1 476.06 ;
      RECT 3.12 478.86 6.84 479.66 ;
      RECT 3.12 479.06 88.1 479.46 ;
      RECT 3.12 482.26 6.84 483.06 ;
      RECT 3.12 482.46 88.1 482.86 ;
      RECT 3.12 485.66 6.84 486.46 ;
      RECT 3.12 485.86 88.1 486.26 ;
      RECT 3.12 489.06 6.84 489.86 ;
      RECT 3.12 489.26 88.1 489.66 ;
      RECT 3.12 492.46 6.84 493.26 ;
      RECT 3.12 492.66 88.1 493.06 ;
      RECT 3.12 495.86 6.84 496.66 ;
      RECT 3.12 496.06 88.1 496.46 ;
      RECT 3.12 499.26 6.84 500.06 ;
      RECT 3.12 499.46 88.1 499.86 ;
      RECT 3.12 502.66 6.84 503.46 ;
      RECT 3.12 502.86 88.1 503.26 ;
      RECT 86.61 510.34 87.41 510.94 ;
      RECT 85.41 510.34 86.21 510.94 ;
      RECT 85.41 510.34 87.41 510.74 ;
      RECT 86.9 7.09 87.22 7.9 ;
      RECT 86.96 7.04 87.16 7.9 ;
      RECT 84.51 67.59 86.61 68.59 ;
      RECT 86.21 6.24 86.61 68.59 ;
      RECT 84.91 37.61 85.51 37.81 ;
      RECT 84.91 28.55 85.11 37.81 ;
      RECT 85.31 28.55 85.51 37.41 ;
      RECT 84.91 28.55 86.61 28.75 ;
      RECT 85.51 28.15 86.61 28.75 ;
      RECT 85.41 6.24 86.71 6.84 ;
      RECT 85.31 38.01 85.51 65.45 ;
      RECT 85.31 38.01 85.91 38.21 ;
      RECT 85.71 30.13 85.91 38.21 ;
      RECT 83.81 27.82 84.21 68.59 ;
      RECT 82.11 65.96 85.91 66.96 ;
      RECT 84.21 6.24 84.95 28.22 ;
      RECT 83.03 6.24 84.95 18.31 ;
      RECT 83.03 6.24 85.01 7.44 ;
      RECT 84.91 38.01 85.11 65.05 ;
      RECT 84.51 38.01 85.11 38.21 ;
      RECT 84.51 30.13 84.71 38.21 ;
      RECT 82.91 38.01 83.11 65.05 ;
      RECT 82.91 38.01 83.51 38.21 ;
      RECT 83.31 30.13 83.51 38.21 ;
      RECT 79.71 67.59 83.51 68.59 ;
      RECT 81.41 28.15 81.81 68.59 ;
      RECT 82.51 37.61 83.11 37.81 ;
      RECT 82.91 28.75 83.11 37.81 ;
      RECT 82.51 28.15 82.71 37.41 ;
      RECT 82.51 28.75 83.11 28.95 ;
      RECT 82.51 38.01 82.71 65.45 ;
      RECT 82.11 38.01 82.71 38.21 ;
      RECT 82.11 30.13 82.31 38.21 ;
      RECT 80.91 6.24 82.31 25.07 ;
      RECT 80.63 6.24 82.61 7.44 ;
      RECT 81.81 510.34 82.61 510.94 ;
      RECT 80.61 510.34 81.41 510.94 ;
      RECT 80.61 510.34 82.61 510.74 ;
      RECT 80.51 38.01 80.71 65.45 ;
      RECT 80.51 38.01 81.11 38.21 ;
      RECT 80.91 30.13 81.11 38.21 ;
      RECT 79.01 27.82 79.41 68.59 ;
      RECT 77.31 65.96 81.11 66.96 ;
      RECT 78.27 6.24 79.01 28.22 ;
      RECT 78.27 6.24 80.21 18.31 ;
      RECT 78.23 6.24 80.21 7.44 ;
      RECT 80.11 37.61 80.71 37.81 ;
      RECT 80.11 28.75 80.31 37.81 ;
      RECT 80.51 28.15 80.71 37.41 ;
      RECT 80.11 28.75 80.71 28.95 ;
      RECT 80.11 38.01 80.31 65.05 ;
      RECT 79.71 38.01 80.31 38.21 ;
      RECT 79.71 30.13 79.91 38.21 ;
      RECT 78.11 38.01 78.31 65.05 ;
      RECT 78.11 38.01 78.71 38.21 ;
      RECT 78.51 30.13 78.71 38.21 ;
      RECT 74.91 67.59 78.71 68.59 ;
      RECT 76.61 6.24 77.01 68.59 ;
      RECT 77.71 37.61 78.31 37.81 ;
      RECT 78.11 28.55 78.31 37.81 ;
      RECT 75.31 37.61 75.91 37.81 ;
      RECT 75.31 28.55 75.51 37.81 ;
      RECT 77.71 28.55 77.91 37.41 ;
      RECT 75.71 28.55 75.91 37.41 ;
      RECT 75.71 28.55 77.01 28.95 ;
      RECT 75.31 28.55 78.31 28.75 ;
      RECT 76.61 28.15 77.71 28.75 ;
      RECT 76.21 9.34 77.01 9.54 ;
      RECT 75.81 6.24 77.81 6.84 ;
      RECT 77.71 38.01 77.91 65.45 ;
      RECT 77.31 38.01 77.91 38.21 ;
      RECT 77.31 30.13 77.51 38.21 ;
      RECT 77.01 510.34 77.81 510.94 ;
      RECT 75.81 510.34 76.61 510.94 ;
      RECT 75.81 510.34 77.81 510.74 ;
      RECT 75.71 38.01 75.91 65.45 ;
      RECT 75.71 38.01 76.31 38.21 ;
      RECT 76.11 30.13 76.31 38.21 ;
      RECT 74.21 27.82 74.61 68.59 ;
      RECT 72.51 65.96 76.31 66.96 ;
      RECT 74.21 27.82 75.35 28.22 ;
      RECT 75.15 7.54 75.35 28.22 ;
      RECT 74.61 7.54 75.35 20.81 ;
      RECT 74.21 6.24 75.01 8.24 ;
      RECT 73.44 6.24 75.41 6.84 ;
      RECT 75.96 25.29 76.16 28.35 ;
      RECT 75.75 25.29 76.16 25.49 ;
      RECT 75.75 21.25 75.95 25.49 ;
      RECT 75.31 38.01 75.51 65.05 ;
      RECT 74.91 38.01 75.51 38.21 ;
      RECT 74.91 30.13 75.11 38.21 ;
      RECT 73.81 27.42 74.01 28.57 ;
      RECT 73.81 27.42 74.95 27.62 ;
      RECT 74.75 21.01 74.95 27.62 ;
      RECT 74.21 21.01 74.95 21.21 ;
      RECT 74.21 18.71 74.41 21.21 ;
      RECT 72.91 37.61 73.51 37.81 ;
      RECT 73.31 27.02 73.51 37.81 ;
      RECT 73.31 27.02 74.55 27.22 ;
      RECT 74.35 21.41 74.55 27.22 ;
      RECT 73.81 21.41 74.55 21.61 ;
      RECT 73.81 12.98 74.01 21.61 ;
      RECT 73.95 21.81 74.15 23.85 ;
      RECT 73.41 21.81 74.15 22.01 ;
      RECT 73.41 20.73 73.61 22.01 ;
      RECT 73.31 38.01 73.51 65.05 ;
      RECT 73.31 38.01 73.91 38.21 ;
      RECT 73.71 30.13 73.91 38.21 ;
      RECT 70.11 67.59 73.91 68.59 ;
      RECT 71.81 26.07 72.21 68.59 ;
      RECT 71.31 26.07 72.21 28.61 ;
      RECT 71.31 26.07 72.71 28.6 ;
      RECT 70.65 26.07 73.37 26.27 ;
      RECT 73.17 24.87 73.37 26.27 ;
      RECT 70.65 24.87 70.85 26.27 ;
      RECT 70.65 24.87 73.37 25.07 ;
      RECT 71.31 14.44 72.71 25.07 ;
      RECT 71.81 6.24 72.21 25.07 ;
      RECT 71.51 6.24 73.01 6.84 ;
      RECT 72.91 38.01 73.11 65.45 ;
      RECT 72.51 38.01 73.11 38.21 ;
      RECT 72.51 30.13 72.71 38.21 ;
      RECT 72.21 510.34 73.01 510.94 ;
      RECT 71.01 510.34 71.81 510.94 ;
      RECT 71.01 510.34 73.01 510.74 ;
      RECT 70.51 37.61 71.11 37.81 ;
      RECT 70.51 27.02 70.71 37.81 ;
      RECT 69.47 27.02 70.71 27.22 ;
      RECT 69.47 21.41 69.67 27.22 ;
      RECT 69.47 21.41 70.21 21.61 ;
      RECT 70.01 19.42 70.21 21.61 ;
      RECT 70.01 19.42 70.81 19.62 ;
      RECT 70.61 13.78 70.81 19.62 ;
      RECT 70.61 13.78 71.61 13.98 ;
      RECT 71.41 8.94 71.61 13.98 ;
      RECT 70.91 38.01 71.11 65.45 ;
      RECT 70.91 38.01 71.51 38.21 ;
      RECT 71.31 30.13 71.51 38.21 ;
      RECT 69.41 27.82 69.81 68.59 ;
      RECT 67.71 65.96 71.51 66.96 ;
      RECT 68.67 27.82 69.81 28.22 ;
      RECT 68.67 7.54 68.87 28.22 ;
      RECT 68.67 16.1 69.41 20.81 ;
      RECT 68.27 14.76 69.01 16.84 ;
      RECT 68.67 7.54 69.41 15.5 ;
      RECT 69.11 6.24 69.91 8.24 ;
      RECT 69.11 6.24 70.11 6.84 ;
      RECT 71.01 8.94 71.21 13.58 ;
      RECT 70.74 8.94 71.21 9.14 ;
      RECT 70.51 38.01 70.71 65.05 ;
      RECT 70.11 38.01 70.71 38.21 ;
      RECT 70.11 30.13 70.31 38.21 ;
      RECT 69.87 21.81 70.07 23.85 ;
      RECT 69.87 21.81 70.61 22.01 ;
      RECT 70.41 20.73 70.61 22.01 ;
      RECT 70.01 27.42 70.21 28.57 ;
      RECT 69.07 27.42 70.21 27.62 ;
      RECT 69.07 21.01 69.27 27.62 ;
      RECT 69.07 21.01 69.81 21.21 ;
      RECT 69.61 15.7 69.81 21.21 ;
      RECT 69.21 15.7 69.81 15.9 ;
      RECT 68.51 38.01 68.71 65.05 ;
      RECT 68.51 38.01 69.11 38.21 ;
      RECT 68.91 30.13 69.11 38.21 ;
      RECT 65.31 67.59 69.11 68.59 ;
      RECT 67.01 6.24 67.41 68.59 ;
      RECT 68.11 37.61 68.71 37.81 ;
      RECT 68.51 28.55 68.71 37.81 ;
      RECT 65.71 37.61 66.31 37.81 ;
      RECT 65.71 28.55 65.91 37.81 ;
      RECT 68.11 28.55 68.31 37.41 ;
      RECT 66.11 28.55 66.31 37.41 ;
      RECT 66.11 28.55 68.31 28.95 ;
      RECT 65.71 28.55 68.71 28.75 ;
      RECT 66.81 6.24 67.61 6.84 ;
      RECT 67.61 9.82 67.81 15.58 ;
      RECT 67.61 9.82 68.31 10.02 ;
      RECT 68.11 7.14 68.31 10.02 ;
      RECT 68.11 38.01 68.31 65.45 ;
      RECT 67.71 38.01 68.31 38.21 ;
      RECT 67.71 30.13 67.91 38.21 ;
      RECT 67.86 25.29 68.06 28.35 ;
      RECT 67.86 25.29 68.27 25.49 ;
      RECT 68.07 21.25 68.27 25.49 ;
      RECT 67.41 510.34 68.21 510.94 ;
      RECT 66.21 510.34 67.01 510.94 ;
      RECT 66.21 510.34 68.21 510.74 ;
      RECT 66.61 9.82 66.81 15.58 ;
      RECT 66.11 9.82 66.81 10.02 ;
      RECT 66.11 7.14 66.31 10.02 ;
      RECT 66.11 38.01 66.31 65.45 ;
      RECT 66.11 38.01 66.71 38.21 ;
      RECT 66.51 30.13 66.71 38.21 ;
      RECT 64.61 27.82 65.01 68.59 ;
      RECT 62.91 65.96 66.71 66.96 ;
      RECT 64.61 27.82 65.75 28.22 ;
      RECT 65.55 7.54 65.75 28.22 ;
      RECT 65.01 16.1 65.75 20.81 ;
      RECT 65.41 14.76 66.15 16.84 ;
      RECT 65.01 7.54 65.75 15.5 ;
      RECT 64.51 6.24 65.31 8.24 ;
      RECT 64.31 6.24 65.31 6.84 ;
      RECT 66.36 25.29 66.56 28.35 ;
      RECT 66.15 25.29 66.56 25.49 ;
      RECT 66.15 21.25 66.35 25.49 ;
      RECT 65.71 38.01 65.91 65.05 ;
      RECT 65.31 38.01 65.91 38.21 ;
      RECT 65.31 30.13 65.51 38.21 ;
      RECT 64.21 27.42 64.41 28.57 ;
      RECT 64.21 27.42 65.35 27.62 ;
      RECT 65.15 21.01 65.35 27.62 ;
      RECT 64.61 21.01 65.35 21.21 ;
      RECT 64.61 15.7 64.81 21.21 ;
      RECT 64.61 15.7 65.21 15.9 ;
      RECT 63.31 37.61 63.91 37.81 ;
      RECT 63.71 27.02 63.91 37.81 ;
      RECT 63.71 27.02 64.95 27.22 ;
      RECT 64.75 21.41 64.95 27.22 ;
      RECT 64.21 21.41 64.95 21.61 ;
      RECT 64.21 19.42 64.41 21.61 ;
      RECT 63.61 19.42 64.41 19.62 ;
      RECT 63.61 13.78 63.81 19.62 ;
      RECT 62.81 13.78 63.81 13.98 ;
      RECT 62.81 8.94 63.01 13.98 ;
      RECT 64.35 21.81 64.55 23.85 ;
      RECT 63.81 21.81 64.55 22.01 ;
      RECT 63.81 20.73 64.01 22.01 ;
      RECT 63.71 38.01 63.91 65.05 ;
      RECT 63.71 38.01 64.31 38.21 ;
      RECT 64.11 30.13 64.31 38.21 ;
      RECT 60.51 67.59 64.31 68.59 ;
      RECT 62.21 26.07 62.61 68.59 ;
      RECT 62.21 26.07 63.11 28.61 ;
      RECT 61.71 26.07 63.11 28.6 ;
      RECT 61.05 26.07 63.77 26.27 ;
      RECT 63.57 24.87 63.77 26.27 ;
      RECT 61.05 24.87 61.25 26.27 ;
      RECT 61.05 24.87 63.77 25.07 ;
      RECT 61.71 14.44 63.11 25.07 ;
      RECT 62.21 6.24 62.61 25.07 ;
      RECT 61.41 6.24 62.91 6.84 ;
      RECT 63.21 8.94 63.41 13.58 ;
      RECT 63.21 8.94 63.68 9.14 ;
      RECT 63.31 38.01 63.51 65.45 ;
      RECT 62.91 38.01 63.51 38.21 ;
      RECT 62.91 30.13 63.11 38.21 ;
      RECT 62.61 510.34 63.41 510.94 ;
      RECT 61.41 510.34 62.21 510.94 ;
      RECT 61.41 510.34 63.41 510.74 ;
      RECT 61.31 38.01 61.51 65.45 ;
      RECT 61.31 38.01 61.91 38.21 ;
      RECT 61.71 30.13 61.91 38.21 ;
      RECT 59.81 27.82 60.21 68.59 ;
      RECT 58.11 65.96 61.91 66.96 ;
      RECT 59.07 27.82 60.21 28.22 ;
      RECT 59.07 7.54 59.27 28.22 ;
      RECT 59.07 7.54 59.81 20.81 ;
      RECT 59.41 6.24 60.21 8.24 ;
      RECT 59.01 6.24 60.98 6.84 ;
      RECT 60.91 37.61 61.51 37.81 ;
      RECT 60.91 27.02 61.11 37.81 ;
      RECT 59.87 27.02 61.11 27.22 ;
      RECT 59.87 21.41 60.07 27.22 ;
      RECT 59.87 21.41 60.61 21.61 ;
      RECT 60.41 12.98 60.61 21.61 ;
      RECT 60.91 38.01 61.11 65.05 ;
      RECT 60.51 38.01 61.11 38.21 ;
      RECT 60.51 30.13 60.71 38.21 ;
      RECT 60.27 21.81 60.47 23.85 ;
      RECT 60.27 21.81 61.01 22.01 ;
      RECT 60.81 20.73 61.01 22.01 ;
      RECT 60.41 27.42 60.61 28.57 ;
      RECT 59.47 27.42 60.61 27.62 ;
      RECT 59.47 21.01 59.67 27.62 ;
      RECT 59.47 21.01 60.21 21.21 ;
      RECT 60.01 18.71 60.21 21.21 ;
      RECT 58.91 38.01 59.11 65.05 ;
      RECT 58.91 38.01 59.51 38.21 ;
      RECT 59.31 30.13 59.51 38.21 ;
      RECT 55.71 67.59 59.51 68.59 ;
      RECT 57.41 6.24 57.81 68.59 ;
      RECT 58.51 37.61 59.11 37.81 ;
      RECT 58.91 28.55 59.11 37.81 ;
      RECT 56.11 37.61 56.71 37.81 ;
      RECT 56.11 28.55 56.31 37.81 ;
      RECT 58.51 28.55 58.71 37.41 ;
      RECT 56.51 28.55 56.71 37.41 ;
      RECT 57.41 28.55 58.71 28.95 ;
      RECT 56.11 28.55 59.11 28.75 ;
      RECT 56.71 28.15 57.81 28.75 ;
      RECT 57.41 9.34 58.21 9.54 ;
      RECT 56.61 6.24 58.61 6.84 ;
      RECT 58.51 38.01 58.71 65.45 ;
      RECT 58.11 38.01 58.71 38.21 ;
      RECT 58.11 30.13 58.31 38.21 ;
      RECT 58.26 25.29 58.46 28.35 ;
      RECT 58.26 25.29 58.67 25.49 ;
      RECT 58.47 21.25 58.67 25.49 ;
      RECT 57.81 510.34 58.61 510.94 ;
      RECT 56.61 510.34 57.41 510.94 ;
      RECT 56.61 510.34 58.61 510.74 ;
      RECT 56.51 38.01 56.71 65.45 ;
      RECT 56.51 38.01 57.11 38.21 ;
      RECT 56.91 30.13 57.11 38.21 ;
      RECT 55.01 27.82 55.41 68.59 ;
      RECT 53.31 65.96 57.11 66.96 ;
      RECT 55.41 6.24 56.15 28.22 ;
      RECT 54.21 6.24 56.15 18.31 ;
      RECT 54.21 6.24 56.19 7.44 ;
      RECT 56.11 38.01 56.31 65.05 ;
      RECT 55.71 38.01 56.31 38.21 ;
      RECT 55.71 30.13 55.91 38.21 ;
      RECT 54.11 38.01 54.31 65.05 ;
      RECT 54.11 38.01 54.71 38.21 ;
      RECT 54.51 30.13 54.71 38.21 ;
      RECT 50.91 67.59 54.71 68.59 ;
      RECT 52.61 28.15 53.01 68.59 ;
      RECT 53.71 37.61 54.31 37.81 ;
      RECT 54.11 28.75 54.31 37.81 ;
      RECT 53.71 28.15 53.91 37.41 ;
      RECT 53.71 28.75 54.31 28.95 ;
      RECT 53.71 38.01 53.91 65.45 ;
      RECT 53.31 38.01 53.91 38.21 ;
      RECT 53.31 30.13 53.51 38.21 ;
      RECT 53.01 510.34 53.81 510.94 ;
      RECT 51.81 510.34 52.61 510.94 ;
      RECT 51.81 510.34 53.81 510.74 ;
      RECT 52.11 6.24 53.51 25.07 ;
      RECT 51.81 6.24 53.79 7.44 ;
      RECT 51.71 38.01 51.91 65.45 ;
      RECT 51.71 38.01 52.31 38.21 ;
      RECT 52.11 30.13 52.31 38.21 ;
      RECT 50.21 27.82 50.61 68.59 ;
      RECT 48.51 65.96 52.31 66.96 ;
      RECT 49.47 6.24 50.21 28.22 ;
      RECT 49.47 6.24 51.39 18.31 ;
      RECT 49.41 6.24 51.39 7.44 ;
      RECT 51.31 37.61 51.91 37.81 ;
      RECT 51.31 28.75 51.51 37.81 ;
      RECT 51.71 28.15 51.91 37.41 ;
      RECT 51.31 28.75 51.91 28.95 ;
      RECT 51.31 38.01 51.51 65.05 ;
      RECT 50.91 38.01 51.51 38.21 ;
      RECT 50.91 30.13 51.11 38.21 ;
      RECT 49.31 38.01 49.51 65.05 ;
      RECT 49.31 38.01 49.91 38.21 ;
      RECT 49.71 30.13 49.91 38.21 ;
      RECT 47.81 67.59 49.91 68.59 ;
      RECT 44.91 67.59 47.01 68.59 ;
      RECT 46.61 6.24 47.01 68.59 ;
      RECT 47.81 6.24 48.21 68.59 ;
      RECT 47.21 7.04 47.61 55.22 ;
      RECT 48.91 37.61 49.51 37.81 ;
      RECT 49.31 28.55 49.51 37.81 ;
      RECT 45.31 37.61 45.91 37.81 ;
      RECT 45.31 28.55 45.51 37.81 ;
      RECT 48.91 28.55 49.11 37.41 ;
      RECT 45.71 28.55 45.91 37.41 ;
      RECT 47.81 28.55 49.51 28.75 ;
      RECT 45.31 28.55 47.01 28.75 ;
      RECT 45.91 28.15 47.01 28.75 ;
      RECT 47.81 28.15 48.91 28.75 ;
      RECT 47.61 6.24 48.21 9.04 ;
      RECT 46.61 6.24 47.21 9.04 ;
      RECT 47.61 6.24 49.01 6.84 ;
      RECT 45.81 6.24 47.21 6.84 ;
      RECT 48.91 38.01 49.11 65.45 ;
      RECT 48.51 38.01 49.11 38.21 ;
      RECT 48.51 30.13 48.71 38.21 ;
      RECT 48.21 510.34 49.01 510.94 ;
      RECT 47.01 510.34 47.81 510.94 ;
      RECT 45.81 510.34 46.61 510.94 ;
      RECT 45.81 510.34 49.01 510.74 ;
      RECT 45.71 38.01 45.91 65.45 ;
      RECT 45.71 38.01 46.31 38.21 ;
      RECT 46.11 30.13 46.31 38.21 ;
      RECT 44.21 27.82 44.61 68.59 ;
      RECT 42.51 65.96 46.31 66.96 ;
      RECT 44.61 6.24 45.35 28.22 ;
      RECT 43.43 6.24 45.35 18.31 ;
      RECT 43.43 6.24 45.41 7.44 ;
      RECT 45.31 38.01 45.51 65.05 ;
      RECT 44.91 38.01 45.51 38.21 ;
      RECT 44.91 30.13 45.11 38.21 ;
      RECT 3.12 508.1 45.19 508.6 ;
      RECT 44.69 506.4 45.19 508.6 ;
      RECT 3.12 506.6 7.71 508.6 ;
      RECT 3.12 507.3 45.19 507.7 ;
      RECT 7.2 506.4 45.19 506.9 ;
      RECT 43.31 38.01 43.51 65.05 ;
      RECT 43.31 38.01 43.91 38.21 ;
      RECT 43.71 30.13 43.91 38.21 ;
      RECT 40.11 67.59 43.91 68.59 ;
      RECT 41.81 28.15 42.21 68.59 ;
      RECT 42.91 37.61 43.51 37.81 ;
      RECT 43.31 28.75 43.51 37.81 ;
      RECT 42.91 28.15 43.11 37.41 ;
      RECT 42.91 28.75 43.51 28.95 ;
      RECT 42.91 38.01 43.11 65.45 ;
      RECT 42.51 38.01 43.11 38.21 ;
      RECT 42.51 30.13 42.71 38.21 ;
      RECT 41.31 6.24 42.71 25.07 ;
      RECT 41.03 6.24 43.01 7.44 ;
      RECT 42.21 510.34 43.01 510.94 ;
      RECT 41.01 510.34 41.81 510.94 ;
      RECT 41.01 510.34 43.01 510.74 ;
      RECT 40.91 38.01 41.11 65.45 ;
      RECT 40.91 38.01 41.51 38.21 ;
      RECT 41.31 30.13 41.51 38.21 ;
      RECT 39.41 27.82 39.81 68.59 ;
      RECT 37.71 65.96 41.51 66.96 ;
      RECT 38.67 6.24 39.41 28.22 ;
      RECT 38.67 6.24 40.61 18.31 ;
      RECT 38.63 6.24 40.61 7.44 ;
      RECT 40.51 37.61 41.11 37.81 ;
      RECT 40.51 28.75 40.71 37.81 ;
      RECT 40.91 28.15 41.11 37.41 ;
      RECT 40.51 28.75 41.11 28.95 ;
      RECT 40.51 38.01 40.71 65.05 ;
      RECT 40.11 38.01 40.71 38.21 ;
      RECT 40.11 30.13 40.31 38.21 ;
      RECT 38.51 38.01 38.71 65.05 ;
      RECT 38.51 38.01 39.11 38.21 ;
      RECT 38.91 30.13 39.11 38.21 ;
      RECT 35.31 67.59 39.11 68.59 ;
      RECT 37.01 6.24 37.41 68.59 ;
      RECT 38.11 37.61 38.71 37.81 ;
      RECT 38.51 28.55 38.71 37.81 ;
      RECT 35.71 37.61 36.31 37.81 ;
      RECT 35.71 28.55 35.91 37.81 ;
      RECT 38.11 28.55 38.31 37.41 ;
      RECT 36.11 28.55 36.31 37.41 ;
      RECT 36.11 28.55 37.41 28.95 ;
      RECT 35.71 28.55 38.71 28.75 ;
      RECT 37.01 28.15 38.11 28.75 ;
      RECT 36.61 9.34 37.41 9.54 ;
      RECT 36.21 6.24 38.21 6.84 ;
      RECT 38.11 38.01 38.31 65.45 ;
      RECT 37.71 38.01 38.31 38.21 ;
      RECT 37.71 30.13 37.91 38.21 ;
      RECT 37.41 510.34 38.21 510.94 ;
      RECT 36.21 510.34 37.01 510.94 ;
      RECT 36.21 510.34 38.21 510.74 ;
      RECT 36.11 38.01 36.31 65.45 ;
      RECT 36.11 38.01 36.71 38.21 ;
      RECT 36.51 30.13 36.71 38.21 ;
      RECT 34.61 27.82 35.01 68.59 ;
      RECT 32.91 65.96 36.71 66.96 ;
      RECT 34.61 27.82 35.75 28.22 ;
      RECT 35.55 7.54 35.75 28.22 ;
      RECT 35.01 7.54 35.75 20.81 ;
      RECT 34.61 6.24 35.41 8.24 ;
      RECT 33.84 6.24 35.81 6.84 ;
      RECT 36.36 25.29 36.56 28.35 ;
      RECT 36.15 25.29 36.56 25.49 ;
      RECT 36.15 21.25 36.35 25.49 ;
      RECT 35.71 38.01 35.91 65.05 ;
      RECT 35.31 38.01 35.91 38.21 ;
      RECT 35.31 30.13 35.51 38.21 ;
      RECT 34.21 27.42 34.41 28.57 ;
      RECT 34.21 27.42 35.35 27.62 ;
      RECT 35.15 21.01 35.35 27.62 ;
      RECT 34.61 21.01 35.35 21.21 ;
      RECT 34.61 18.71 34.81 21.21 ;
      RECT 33.31 37.61 33.91 37.81 ;
      RECT 33.71 27.02 33.91 37.81 ;
      RECT 33.71 27.02 34.95 27.22 ;
      RECT 34.75 21.41 34.95 27.22 ;
      RECT 34.21 21.41 34.95 21.61 ;
      RECT 34.21 12.98 34.41 21.61 ;
      RECT 34.35 21.81 34.55 23.85 ;
      RECT 33.81 21.81 34.55 22.01 ;
      RECT 33.81 20.73 34.01 22.01 ;
      RECT 33.71 38.01 33.91 65.05 ;
      RECT 33.71 38.01 34.31 38.21 ;
      RECT 34.11 30.13 34.31 38.21 ;
      RECT 30.51 67.59 34.31 68.59 ;
      RECT 32.21 26.07 32.61 68.59 ;
      RECT 31.71 26.07 32.61 28.61 ;
      RECT 31.71 26.07 33.11 28.6 ;
      RECT 31.05 26.07 33.77 26.27 ;
      RECT 33.57 24.87 33.77 26.27 ;
      RECT 31.05 24.87 31.25 26.27 ;
      RECT 31.05 24.87 33.77 25.07 ;
      RECT 31.71 14.44 33.11 25.07 ;
      RECT 32.21 6.24 32.61 25.07 ;
      RECT 31.91 6.24 33.41 6.84 ;
      RECT 33.31 38.01 33.51 65.45 ;
      RECT 32.91 38.01 33.51 38.21 ;
      RECT 32.91 30.13 33.11 38.21 ;
      RECT 32.61 510.34 33.41 510.94 ;
      RECT 31.41 510.34 32.21 510.94 ;
      RECT 31.41 510.34 33.41 510.74 ;
      RECT 30.91 37.61 31.51 37.81 ;
      RECT 30.91 27.02 31.11 37.81 ;
      RECT 29.87 27.02 31.11 27.22 ;
      RECT 29.87 21.41 30.07 27.22 ;
      RECT 29.87 21.41 30.61 21.61 ;
      RECT 30.41 19.42 30.61 21.61 ;
      RECT 30.41 19.42 31.21 19.62 ;
      RECT 31.01 13.78 31.21 19.62 ;
      RECT 31.01 13.78 32.01 13.98 ;
      RECT 31.81 8.94 32.01 13.98 ;
      RECT 31.31 38.01 31.51 65.45 ;
      RECT 31.31 38.01 31.91 38.21 ;
      RECT 31.71 30.13 31.91 38.21 ;
      RECT 29.81 27.82 30.21 68.59 ;
      RECT 28.11 65.96 31.91 66.96 ;
      RECT 29.07 27.82 30.21 28.22 ;
      RECT 29.07 7.54 29.27 28.22 ;
      RECT 29.07 16.1 29.81 20.81 ;
      RECT 28.67 14.76 29.41 16.84 ;
      RECT 29.07 7.54 29.81 15.5 ;
      RECT 29.51 6.24 30.31 8.24 ;
      RECT 29.51 6.24 30.51 6.84 ;
      RECT 31.41 8.94 31.61 13.58 ;
      RECT 31.14 8.94 31.61 9.14 ;
      RECT 30.91 38.01 31.11 65.05 ;
      RECT 30.51 38.01 31.11 38.21 ;
      RECT 30.51 30.13 30.71 38.21 ;
      RECT 30.27 21.81 30.47 23.85 ;
      RECT 30.27 21.81 31.01 22.01 ;
      RECT 30.81 20.73 31.01 22.01 ;
      RECT 30.41 27.42 30.61 28.57 ;
      RECT 29.47 27.42 30.61 27.62 ;
      RECT 29.47 21.01 29.67 27.62 ;
      RECT 29.47 21.01 30.21 21.21 ;
      RECT 30.01 15.7 30.21 21.21 ;
      RECT 29.61 15.7 30.21 15.9 ;
      RECT 28.91 38.01 29.11 65.05 ;
      RECT 28.91 38.01 29.51 38.21 ;
      RECT 29.31 30.13 29.51 38.21 ;
      RECT 25.71 67.59 29.51 68.59 ;
      RECT 27.41 6.24 27.81 68.59 ;
      RECT 28.51 37.61 29.11 37.81 ;
      RECT 28.91 28.55 29.11 37.81 ;
      RECT 26.11 37.61 26.71 37.81 ;
      RECT 26.11 28.55 26.31 37.81 ;
      RECT 28.51 28.55 28.71 37.41 ;
      RECT 26.51 28.55 26.71 37.41 ;
      RECT 26.51 28.55 28.71 28.95 ;
      RECT 26.11 28.55 29.11 28.75 ;
      RECT 27.21 6.24 28.01 6.84 ;
      RECT 28.01 9.82 28.21 15.58 ;
      RECT 28.01 9.82 28.71 10.02 ;
      RECT 28.51 7.14 28.71 10.02 ;
      RECT 28.51 38.01 28.71 65.45 ;
      RECT 28.11 38.01 28.71 38.21 ;
      RECT 28.11 30.13 28.31 38.21 ;
      RECT 28.26 25.29 28.46 28.35 ;
      RECT 28.26 25.29 28.67 25.49 ;
      RECT 28.47 21.25 28.67 25.49 ;
      RECT 27.81 510.34 28.61 510.94 ;
      RECT 26.61 510.34 27.41 510.94 ;
      RECT 26.61 510.34 28.61 510.74 ;
      RECT 27.01 9.82 27.21 15.58 ;
      RECT 26.51 9.82 27.21 10.02 ;
      RECT 26.51 7.14 26.71 10.02 ;
      RECT 26.51 38.01 26.71 65.45 ;
      RECT 26.51 38.01 27.11 38.21 ;
      RECT 26.91 30.13 27.11 38.21 ;
      RECT 25.01 27.82 25.41 68.59 ;
      RECT 23.31 65.96 27.11 66.96 ;
      RECT 25.01 27.82 26.15 28.22 ;
      RECT 25.95 7.54 26.15 28.22 ;
      RECT 25.41 16.1 26.15 20.81 ;
      RECT 25.81 14.76 26.55 16.84 ;
      RECT 25.41 7.54 26.15 15.5 ;
      RECT 24.91 6.24 25.71 8.24 ;
      RECT 24.71 6.24 25.71 6.84 ;
      RECT 26.76 25.29 26.96 28.35 ;
      RECT 26.55 25.29 26.96 25.49 ;
      RECT 26.55 21.25 26.75 25.49 ;
      RECT 26.11 38.01 26.31 65.05 ;
      RECT 25.71 38.01 26.31 38.21 ;
      RECT 25.71 30.13 25.91 38.21 ;
      RECT 24.61 27.42 24.81 28.57 ;
      RECT 24.61 27.42 25.75 27.62 ;
      RECT 25.55 21.01 25.75 27.62 ;
      RECT 25.01 21.01 25.75 21.21 ;
      RECT 25.01 15.7 25.21 21.21 ;
      RECT 25.01 15.7 25.61 15.9 ;
      RECT 23.71 37.61 24.31 37.81 ;
      RECT 24.11 27.02 24.31 37.81 ;
      RECT 24.11 27.02 25.35 27.22 ;
      RECT 25.15 21.41 25.35 27.22 ;
      RECT 24.61 21.41 25.35 21.61 ;
      RECT 24.61 19.42 24.81 21.61 ;
      RECT 24.01 19.42 24.81 19.62 ;
      RECT 24.01 13.78 24.21 19.62 ;
      RECT 23.21 13.78 24.21 13.98 ;
      RECT 23.21 8.94 23.41 13.98 ;
      RECT 24.75 21.81 24.95 23.85 ;
      RECT 24.21 21.81 24.95 22.01 ;
      RECT 24.21 20.73 24.41 22.01 ;
      RECT 24.11 38.01 24.31 65.05 ;
      RECT 24.11 38.01 24.71 38.21 ;
      RECT 24.51 30.13 24.71 38.21 ;
      RECT 20.91 67.59 24.71 68.59 ;
      RECT 22.61 26.07 23.01 68.59 ;
      RECT 22.61 26.07 23.51 28.61 ;
      RECT 22.11 26.07 23.51 28.6 ;
      RECT 21.45 26.07 24.17 26.27 ;
      RECT 23.97 24.87 24.17 26.27 ;
      RECT 21.45 24.87 21.65 26.27 ;
      RECT 21.45 24.87 24.17 25.07 ;
      RECT 22.11 14.44 23.51 25.07 ;
      RECT 22.61 6.24 23.01 25.07 ;
      RECT 21.81 6.24 23.31 6.84 ;
      RECT 23.61 8.94 23.81 13.58 ;
      RECT 23.61 8.94 24.08 9.14 ;
      RECT 23.71 38.01 23.91 65.45 ;
      RECT 23.31 38.01 23.91 38.21 ;
      RECT 23.31 30.13 23.51 38.21 ;
      RECT 23.01 510.34 23.81 510.94 ;
      RECT 21.81 510.34 22.61 510.94 ;
      RECT 21.81 510.34 23.81 510.74 ;
      RECT 21.71 38.01 21.91 65.45 ;
      RECT 21.71 38.01 22.31 38.21 ;
      RECT 22.11 30.13 22.31 38.21 ;
      RECT 20.21 27.82 20.61 68.59 ;
      RECT 18.51 65.96 22.31 66.96 ;
      RECT 19.47 27.82 20.61 28.22 ;
      RECT 19.47 7.54 19.67 28.22 ;
      RECT 19.47 7.54 20.21 20.81 ;
      RECT 19.81 6.24 20.61 8.24 ;
      RECT 19.81 6.24 21.41 6.84 ;
      RECT 21.31 37.61 21.91 37.81 ;
      RECT 21.31 27.02 21.51 37.81 ;
      RECT 20.27 27.02 21.51 27.22 ;
      RECT 20.27 21.41 20.47 27.22 ;
      RECT 20.27 21.41 21.01 21.61 ;
      RECT 20.81 12.98 21.01 21.61 ;
      RECT 21.31 38.01 21.51 65.05 ;
      RECT 20.91 38.01 21.51 38.21 ;
      RECT 20.91 30.13 21.11 38.21 ;
      RECT 20.67 21.81 20.87 23.85 ;
      RECT 20.67 21.81 21.41 22.01 ;
      RECT 21.21 20.73 21.41 22.01 ;
      RECT 20.81 27.42 21.01 28.57 ;
      RECT 19.87 27.42 21.01 27.62 ;
      RECT 19.87 21.01 20.07 27.62 ;
      RECT 19.87 21.01 20.61 21.21 ;
      RECT 20.41 18.71 20.61 21.21 ;
      RECT 19.31 38.01 19.51 65.05 ;
      RECT 19.31 38.01 19.91 38.21 ;
      RECT 19.71 30.13 19.91 38.21 ;
      RECT 16.11 67.59 19.91 68.59 ;
      RECT 17.81 6.24 18.21 68.59 ;
      RECT 18.91 37.61 19.51 37.81 ;
      RECT 19.31 28.55 19.51 37.81 ;
      RECT 16.51 37.61 17.11 37.81 ;
      RECT 16.51 28.55 16.71 37.81 ;
      RECT 18.91 28.55 19.11 37.41 ;
      RECT 16.91 28.55 17.11 37.41 ;
      RECT 17.81 28.55 19.11 28.95 ;
      RECT 16.51 28.55 19.51 28.75 ;
      RECT 17.11 28.15 18.21 28.75 ;
      RECT 17.81 9.34 18.61 9.54 ;
      RECT 17.01 6.24 18.41 6.84 ;
      RECT 19.01 6.24 19.21 9.14 ;
      RECT 18.81 6.24 19.41 6.84 ;
      RECT 18.91 38.01 19.11 65.45 ;
      RECT 18.51 38.01 19.11 38.21 ;
      RECT 18.51 30.13 18.71 38.21 ;
      RECT 18.66 25.29 18.86 28.35 ;
      RECT 18.66 25.29 19.07 25.49 ;
      RECT 18.87 21.25 19.07 25.49 ;
      RECT 18.21 510.34 19.01 510.94 ;
      RECT 17.01 510.34 17.81 510.94 ;
      RECT 17.01 510.34 19.01 510.74 ;
      RECT 16.91 38.01 17.11 65.45 ;
      RECT 16.91 38.01 17.51 38.21 ;
      RECT 17.31 30.13 17.51 38.21 ;
      RECT 15.41 27.82 15.81 68.59 ;
      RECT 13.71 65.96 17.51 66.96 ;
      RECT 15.81 6.24 16.55 28.22 ;
      RECT 14.61 6.24 16.55 18.31 ;
      RECT 14.61 6.24 16.59 7.44 ;
      RECT 16.51 38.01 16.71 65.05 ;
      RECT 16.11 38.01 16.71 38.21 ;
      RECT 16.11 30.13 16.31 38.21 ;
      RECT 14.51 38.01 14.71 65.05 ;
      RECT 14.51 38.01 15.11 38.21 ;
      RECT 14.91 30.13 15.11 38.21 ;
      RECT 11.31 67.59 15.11 68.59 ;
      RECT 13.01 28.15 13.41 68.59 ;
      RECT 14.11 37.61 14.71 37.81 ;
      RECT 14.51 28.75 14.71 37.81 ;
      RECT 14.11 28.15 14.31 37.41 ;
      RECT 14.11 28.75 14.71 28.95 ;
      RECT 14.11 38.01 14.31 65.45 ;
      RECT 13.71 38.01 14.31 38.21 ;
      RECT 13.71 30.13 13.91 38.21 ;
      RECT 13.41 510.34 14.21 510.94 ;
      RECT 12.21 510.34 13.01 510.94 ;
      RECT 12.21 510.34 14.21 510.74 ;
      RECT 12.51 6.24 13.91 25.07 ;
      RECT 12.21 6.24 14.19 7.44 ;
      RECT 12.11 38.01 12.31 65.45 ;
      RECT 12.11 38.01 12.71 38.21 ;
      RECT 12.51 30.13 12.71 38.21 ;
      RECT 10.61 27.82 11.01 68.59 ;
      RECT 8.91 65.96 12.71 66.96 ;
      RECT 9.87 6.24 10.61 28.22 ;
      RECT 9.87 6.24 11.79 18.31 ;
      RECT 9.81 6.24 11.79 7.44 ;
      RECT 11.71 37.61 12.31 37.81 ;
      RECT 11.71 28.75 11.91 37.81 ;
      RECT 12.11 28.15 12.31 37.41 ;
      RECT 11.71 28.75 12.31 28.95 ;
      RECT 11.71 38.01 11.91 65.05 ;
      RECT 11.31 38.01 11.91 38.21 ;
      RECT 11.31 30.13 11.51 38.21 ;
      RECT 9.71 38.01 9.91 65.05 ;
      RECT 9.71 38.01 10.31 38.21 ;
      RECT 10.11 30.13 10.31 38.21 ;
      RECT 7.21 67.59 10.31 68.59 ;
      RECT 8.21 6.24 8.61 68.59 ;
      RECT 7.41 6.24 7.81 68.59 ;
      RECT 3.12 54.22 7.81 55.22 ;
      RECT 3.12 41.29 7.81 42.29 ;
      RECT 3.12 39.44 7.81 40.44 ;
      RECT 9.31 37.61 9.91 37.81 ;
      RECT 9.71 28.55 9.91 37.81 ;
      RECT 9.31 28.55 9.51 37.41 ;
      RECT 3.12 32.98 7.81 33.98 ;
      RECT 3.12 31.13 7.81 32.13 ;
      RECT 8.21 28.55 9.91 28.75 ;
      RECT 8.21 28.15 9.31 28.75 ;
      RECT 3.12 21.41 7.81 22.21 ;
      RECT 3.12 12.64 7.81 13.74 ;
      RECT 7.41 6.24 9.41 6.84 ;
      RECT 9.31 38.01 9.51 65.45 ;
      RECT 8.91 38.01 9.51 38.21 ;
      RECT 8.91 30.13 9.11 38.21 ;
      RECT 8.61 510.34 9.41 510.94 ;
      RECT 7.41 510.34 8.21 510.94 ;
      RECT 7.21 510.34 9.41 510.74 ;
      RECT 233.76 7.94 240.6 9.14 ;
      RECT 233.76 17.26 240.6 18.46 ;
      RECT 233.76 25.81 240.6 27.81 ;
      RECT 233.76 35.91 240.6 36.91 ;
      RECT 233.76 50.24 240.6 51.24 ;
      RECT 233.76 57.02 240.6 58.02 ;
      RECT 233.76 60.6 240.6 61.6 ;
      RECT 233.76 62.45 240.6 63.45 ;
      RECT 0 515.18 240.6 517.18 ;
      RECT 2.36 0 238.24 2 ;
      RECT 3.12 512.06 237.48 514.06 ;
      RECT 5.48 3.12 235.12 5.12 ;
      RECT 149.73 70.16 233.4 70.66 ;
      RECT 149.73 71.86 233.4 72.36 ;
      RECT 149.73 73.56 233.4 74.06 ;
      RECT 149.73 75.26 233.4 75.76 ;
      RECT 149.73 76.96 233.4 77.46 ;
      RECT 149.73 78.66 233.4 79.16 ;
      RECT 149.73 80.36 233.4 80.86 ;
      RECT 149.73 82.06 233.4 82.56 ;
      RECT 149.73 83.76 233.4 84.26 ;
      RECT 149.73 85.46 233.4 85.96 ;
      RECT 149.73 87.16 233.4 87.66 ;
      RECT 149.73 88.86 233.4 89.36 ;
      RECT 149.73 90.56 233.4 91.06 ;
      RECT 149.73 92.26 233.4 92.76 ;
      RECT 149.73 93.96 233.4 94.46 ;
      RECT 149.73 95.66 233.4 96.16 ;
      RECT 149.73 97.36 233.4 97.86 ;
      RECT 149.73 99.06 233.4 99.56 ;
      RECT 149.73 100.76 233.4 101.26 ;
      RECT 149.73 102.46 233.4 102.96 ;
      RECT 149.73 104.16 233.4 104.66 ;
      RECT 149.73 105.86 233.4 106.36 ;
      RECT 149.73 107.56 233.4 108.06 ;
      RECT 149.73 109.26 233.4 109.76 ;
      RECT 149.73 110.96 233.4 111.46 ;
      RECT 149.73 112.66 233.4 113.16 ;
      RECT 149.73 114.36 233.4 114.86 ;
      RECT 149.73 116.06 233.4 116.56 ;
      RECT 149.73 117.76 233.4 118.26 ;
      RECT 149.73 119.46 233.4 119.96 ;
      RECT 149.73 121.16 233.4 121.66 ;
      RECT 149.73 122.86 233.4 123.36 ;
      RECT 149.73 124.56 233.4 125.06 ;
      RECT 149.73 126.26 233.4 126.76 ;
      RECT 149.73 127.96 233.4 128.46 ;
      RECT 149.73 129.66 233.4 130.16 ;
      RECT 149.73 131.36 233.4 131.86 ;
      RECT 149.73 133.06 233.4 133.56 ;
      RECT 149.73 134.76 233.4 135.26 ;
      RECT 149.73 136.46 233.4 136.96 ;
      RECT 149.73 138.16 233.4 138.66 ;
      RECT 149.73 139.86 233.4 140.36 ;
      RECT 149.73 141.56 233.4 142.06 ;
      RECT 149.73 143.26 233.4 143.76 ;
      RECT 149.73 144.96 233.4 145.46 ;
      RECT 149.73 146.66 233.4 147.16 ;
      RECT 149.73 148.36 233.4 148.86 ;
      RECT 149.73 150.06 233.4 150.56 ;
      RECT 149.73 151.76 233.4 152.26 ;
      RECT 149.73 153.46 233.4 153.96 ;
      RECT 149.73 155.16 233.4 155.66 ;
      RECT 149.73 156.86 233.4 157.36 ;
      RECT 149.73 158.56 233.4 159.06 ;
      RECT 149.73 160.26 233.4 160.76 ;
      RECT 149.73 161.96 233.4 162.46 ;
      RECT 149.73 163.66 233.4 164.16 ;
      RECT 149.73 165.36 233.4 165.86 ;
      RECT 149.73 167.06 233.4 167.56 ;
      RECT 149.73 168.76 233.4 169.26 ;
      RECT 149.73 170.46 233.4 170.96 ;
      RECT 149.73 172.16 233.4 172.66 ;
      RECT 149.73 173.86 233.4 174.36 ;
      RECT 149.73 175.56 233.4 176.06 ;
      RECT 149.73 177.26 233.4 177.76 ;
      RECT 149.73 178.96 233.4 179.46 ;
      RECT 149.73 180.66 233.4 181.16 ;
      RECT 149.73 182.36 233.4 182.86 ;
      RECT 149.73 184.06 233.4 184.56 ;
      RECT 149.73 185.76 233.4 186.26 ;
      RECT 149.73 187.46 233.4 187.96 ;
      RECT 149.73 189.16 233.4 189.66 ;
      RECT 149.73 190.86 233.4 191.36 ;
      RECT 149.73 192.56 233.4 193.06 ;
      RECT 149.73 194.26 233.4 194.76 ;
      RECT 149.73 195.96 233.4 196.46 ;
      RECT 149.73 197.66 233.4 198.16 ;
      RECT 149.73 199.36 233.4 199.86 ;
      RECT 149.73 201.06 233.4 201.56 ;
      RECT 149.73 202.76 233.4 203.26 ;
      RECT 149.73 204.46 233.4 204.96 ;
      RECT 149.73 206.16 233.4 206.66 ;
      RECT 149.73 207.86 233.4 208.36 ;
      RECT 149.73 209.56 233.4 210.06 ;
      RECT 149.73 211.26 233.4 211.76 ;
      RECT 149.73 212.96 233.4 213.46 ;
      RECT 149.73 214.66 233.4 215.16 ;
      RECT 149.73 216.36 233.4 216.86 ;
      RECT 149.73 218.06 233.4 218.56 ;
      RECT 149.73 219.76 233.4 220.26 ;
      RECT 149.73 221.46 233.4 221.96 ;
      RECT 149.73 223.16 233.4 223.66 ;
      RECT 149.73 224.86 233.4 225.36 ;
      RECT 149.73 226.56 233.4 227.06 ;
      RECT 149.73 228.26 233.4 228.76 ;
      RECT 149.73 229.96 233.4 230.46 ;
      RECT 149.73 231.66 233.4 232.16 ;
      RECT 149.73 233.36 233.4 233.86 ;
      RECT 149.73 235.06 233.4 235.56 ;
      RECT 149.73 236.76 233.4 237.26 ;
      RECT 149.73 238.46 233.4 238.96 ;
      RECT 149.73 240.16 233.4 240.66 ;
      RECT 149.73 241.86 233.4 242.36 ;
      RECT 149.73 243.56 233.4 244.06 ;
      RECT 149.73 245.26 233.4 245.76 ;
      RECT 149.73 246.96 233.4 247.46 ;
      RECT 149.73 248.66 233.4 249.16 ;
      RECT 149.73 250.36 233.4 250.86 ;
      RECT 149.73 252.06 233.4 252.56 ;
      RECT 149.73 253.76 233.4 254.26 ;
      RECT 149.73 255.46 233.4 255.96 ;
      RECT 149.73 257.16 233.4 257.66 ;
      RECT 149.73 258.86 233.4 259.36 ;
      RECT 149.73 260.56 233.4 261.06 ;
      RECT 149.73 262.26 233.4 262.76 ;
      RECT 149.73 263.96 233.4 264.46 ;
      RECT 149.73 265.66 233.4 266.16 ;
      RECT 149.73 267.36 233.4 267.86 ;
      RECT 149.73 269.06 233.4 269.56 ;
      RECT 149.73 270.76 233.4 271.26 ;
      RECT 149.73 272.46 233.4 272.96 ;
      RECT 149.73 274.16 233.4 274.66 ;
      RECT 149.73 275.86 233.4 276.36 ;
      RECT 149.73 277.56 233.4 278.06 ;
      RECT 149.73 279.26 233.4 279.76 ;
      RECT 149.73 280.96 233.4 281.46 ;
      RECT 149.73 282.66 233.4 283.16 ;
      RECT 149.73 284.36 233.4 284.86 ;
      RECT 149.73 286.06 233.4 286.56 ;
      RECT 149.73 287.76 233.4 288.26 ;
      RECT 149.73 289.46 233.4 289.96 ;
      RECT 149.73 291.16 233.4 291.66 ;
      RECT 149.73 292.86 233.4 293.36 ;
      RECT 149.73 294.56 233.4 295.06 ;
      RECT 149.73 296.26 233.4 296.76 ;
      RECT 149.73 297.96 233.4 298.46 ;
      RECT 149.73 299.66 233.4 300.16 ;
      RECT 149.73 301.36 233.4 301.86 ;
      RECT 149.73 303.06 233.4 303.56 ;
      RECT 149.73 304.76 233.4 305.26 ;
      RECT 149.73 306.46 233.4 306.96 ;
      RECT 149.73 308.16 233.4 308.66 ;
      RECT 149.73 309.86 233.4 310.36 ;
      RECT 149.73 311.56 233.4 312.06 ;
      RECT 149.73 313.26 233.4 313.76 ;
      RECT 149.73 314.96 233.4 315.46 ;
      RECT 149.73 316.66 233.4 317.16 ;
      RECT 149.73 318.36 233.4 318.86 ;
      RECT 149.73 320.06 233.4 320.56 ;
      RECT 149.73 321.76 233.4 322.26 ;
      RECT 149.73 323.46 233.4 323.96 ;
      RECT 149.73 325.16 233.4 325.66 ;
      RECT 149.73 326.86 233.4 327.36 ;
      RECT 149.73 328.56 233.4 329.06 ;
      RECT 149.73 330.26 233.4 330.76 ;
      RECT 149.73 331.96 233.4 332.46 ;
      RECT 149.73 333.66 233.4 334.16 ;
      RECT 149.73 335.36 233.4 335.86 ;
      RECT 149.73 337.06 233.4 337.56 ;
      RECT 149.73 338.76 233.4 339.26 ;
      RECT 149.73 340.46 233.4 340.96 ;
      RECT 149.73 342.16 233.4 342.66 ;
      RECT 149.73 343.86 233.4 344.36 ;
      RECT 149.73 345.56 233.4 346.06 ;
      RECT 149.73 347.26 233.4 347.76 ;
      RECT 149.73 348.96 233.4 349.46 ;
      RECT 149.73 350.66 233.4 351.16 ;
      RECT 149.73 352.36 233.4 352.86 ;
      RECT 149.73 354.06 233.4 354.56 ;
      RECT 149.73 355.76 233.4 356.26 ;
      RECT 149.73 357.46 233.4 357.96 ;
      RECT 149.73 359.16 233.4 359.66 ;
      RECT 149.73 360.86 233.4 361.36 ;
      RECT 149.73 362.56 233.4 363.06 ;
      RECT 149.73 364.26 233.4 364.76 ;
      RECT 149.73 365.96 233.4 366.46 ;
      RECT 149.73 367.66 233.4 368.16 ;
      RECT 149.73 369.36 233.4 369.86 ;
      RECT 149.73 371.06 233.4 371.56 ;
      RECT 149.73 372.76 233.4 373.26 ;
      RECT 149.73 374.46 233.4 374.96 ;
      RECT 149.73 376.16 233.4 376.66 ;
      RECT 149.73 377.86 233.4 378.36 ;
      RECT 149.73 379.56 233.4 380.06 ;
      RECT 149.73 381.26 233.4 381.76 ;
      RECT 149.73 382.96 233.4 383.46 ;
      RECT 149.73 384.66 233.4 385.16 ;
      RECT 149.73 386.36 233.4 386.86 ;
      RECT 149.73 388.06 233.4 388.56 ;
      RECT 149.73 389.76 233.4 390.26 ;
      RECT 149.73 391.46 233.4 391.96 ;
      RECT 149.73 393.16 233.4 393.66 ;
      RECT 149.73 394.86 233.4 395.36 ;
      RECT 149.73 396.56 233.4 397.06 ;
      RECT 149.73 398.26 233.4 398.76 ;
      RECT 149.73 399.96 233.4 400.46 ;
      RECT 149.73 401.66 233.4 402.16 ;
      RECT 149.73 403.36 233.4 403.86 ;
      RECT 149.73 405.06 233.4 405.56 ;
      RECT 149.73 406.76 233.4 407.26 ;
      RECT 149.73 408.46 233.4 408.96 ;
      RECT 149.73 410.16 233.4 410.66 ;
      RECT 149.73 411.86 233.4 412.36 ;
      RECT 149.73 413.56 233.4 414.06 ;
      RECT 149.73 415.26 233.4 415.76 ;
      RECT 149.73 416.96 233.4 417.46 ;
      RECT 149.73 418.66 233.4 419.16 ;
      RECT 149.73 420.36 233.4 420.86 ;
      RECT 149.73 422.06 233.4 422.56 ;
      RECT 149.73 423.76 233.4 424.26 ;
      RECT 149.73 425.46 233.4 425.96 ;
      RECT 149.73 427.16 233.4 427.66 ;
      RECT 149.73 428.86 233.4 429.36 ;
      RECT 149.73 430.56 233.4 431.06 ;
      RECT 149.73 432.26 233.4 432.76 ;
      RECT 149.73 433.96 233.4 434.46 ;
      RECT 149.73 435.66 233.4 436.16 ;
      RECT 149.73 437.36 233.4 437.86 ;
      RECT 149.73 439.06 233.4 439.56 ;
      RECT 149.73 440.76 233.4 441.26 ;
      RECT 149.73 442.46 233.4 442.96 ;
      RECT 149.73 444.16 233.4 444.66 ;
      RECT 149.73 445.86 233.4 446.36 ;
      RECT 149.73 447.56 233.4 448.06 ;
      RECT 149.73 449.26 233.4 449.76 ;
      RECT 149.73 450.96 233.4 451.46 ;
      RECT 149.73 452.66 233.4 453.16 ;
      RECT 149.73 454.36 233.4 454.86 ;
      RECT 149.73 456.06 233.4 456.56 ;
      RECT 149.73 457.76 233.4 458.26 ;
      RECT 149.73 459.46 233.4 459.96 ;
      RECT 149.73 461.16 233.4 461.66 ;
      RECT 149.73 462.86 233.4 463.36 ;
      RECT 149.73 464.56 233.4 465.06 ;
      RECT 149.73 466.26 233.4 466.76 ;
      RECT 149.73 467.96 233.4 468.46 ;
      RECT 149.73 469.66 233.4 470.16 ;
      RECT 149.73 471.36 233.4 471.86 ;
      RECT 149.73 473.06 233.4 473.56 ;
      RECT 149.73 474.76 233.4 475.26 ;
      RECT 149.73 476.46 233.4 476.96 ;
      RECT 149.73 478.16 233.4 478.66 ;
      RECT 149.73 479.86 233.4 480.36 ;
      RECT 149.73 481.56 233.4 482.06 ;
      RECT 149.73 483.26 233.4 483.76 ;
      RECT 149.73 484.96 233.4 485.46 ;
      RECT 149.73 486.66 233.4 487.16 ;
      RECT 149.73 488.36 233.4 488.86 ;
      RECT 149.73 490.06 233.4 490.56 ;
      RECT 149.73 491.76 233.4 492.26 ;
      RECT 149.73 493.46 233.4 493.96 ;
      RECT 149.73 495.16 233.4 495.66 ;
      RECT 149.73 496.86 233.4 497.36 ;
      RECT 149.73 498.56 233.4 499.06 ;
      RECT 149.73 500.26 233.4 500.76 ;
      RECT 149.73 501.96 233.4 502.46 ;
      RECT 149.73 503.66 233.4 504.16 ;
      RECT 231.49 38.41 231.69 65.45 ;
      RECT 230.29 38.41 230.49 65.45 ;
      RECT 229.09 38.41 229.29 65.45 ;
      RECT 227.89 38.41 228.09 65.45 ;
      RECT 226.69 38.41 226.89 65.45 ;
      RECT 225.49 38.41 225.69 65.45 ;
      RECT 224.29 38.41 224.49 65.45 ;
      RECT 223.09 38.41 223.29 65.45 ;
      RECT 221.99 13.78 222.19 24.54 ;
      RECT 221.89 38.41 222.09 65.45 ;
      RECT 221.39 7.04 221.59 9.14 ;
      RECT 220.69 38.41 220.89 65.45 ;
      RECT 219.75 8.84 219.95 9.44 ;
      RECT 219.49 38.41 219.69 65.45 ;
      RECT 219.33 22.31 219.53 24.62 ;
      RECT 218.98 15.39 219.18 16.47 ;
      RECT 218.69 27.45 218.89 37.41 ;
      RECT 216.83 25.27 218.75 25.47 ;
      RECT 216.83 25.67 218.75 25.87 ;
      RECT 218.29 38.41 218.49 65.45 ;
      RECT 217.09 38.41 217.29 65.45 ;
      RECT 216.69 27.45 216.89 37.41 ;
      RECT 216.05 22.31 216.25 24.62 ;
      RECT 215.89 38.41 216.09 65.45 ;
      RECT 214.69 38.41 214.89 65.45 ;
      RECT 213.49 38.41 213.69 65.45 ;
      RECT 213.39 16.5 213.59 24.54 ;
      RECT 212.39 16.5 212.59 24.54 ;
      RECT 212.29 38.41 212.49 65.45 ;
      RECT 211.09 38.41 211.29 65.45 ;
      RECT 209.89 38.41 210.09 65.45 ;
      RECT 209.73 22.31 209.93 24.62 ;
      RECT 209.09 27.45 209.29 37.41 ;
      RECT 207.23 25.27 209.15 25.47 ;
      RECT 207.23 25.67 209.15 25.87 ;
      RECT 208.69 38.41 208.89 65.45 ;
      RECT 207.49 38.41 207.69 65.45 ;
      RECT 207.09 27.45 207.29 37.41 ;
      RECT 206.8 15.39 207 16.47 ;
      RECT 206.45 22.31 206.65 24.62 ;
      RECT 206.29 38.41 206.49 65.45 ;
      RECT 206.03 8.84 206.23 9.44 ;
      RECT 205.09 38.41 205.29 65.45 ;
      RECT 204.39 7.04 204.59 9.14 ;
      RECT 203.89 38.41 204.09 65.45 ;
      RECT 203.79 13.78 203.99 24.54 ;
      RECT 202.69 38.41 202.89 65.45 ;
      RECT 201.49 38.41 201.69 65.45 ;
      RECT 200.29 38.41 200.49 65.45 ;
      RECT 199.09 38.41 199.29 65.45 ;
      RECT 197.89 38.41 198.09 65.45 ;
      RECT 196.69 38.41 196.89 65.45 ;
      RECT 195.49 38.41 195.69 65.45 ;
      RECT 194.29 38.41 194.49 65.45 ;
      RECT 193.09 57.02 193.29 63.45 ;
      RECT 191.89 38.41 192.09 65.45 ;
      RECT 190.69 38.41 190.89 65.45 ;
      RECT 189.49 38.41 189.69 65.45 ;
      RECT 188.29 38.41 188.49 65.45 ;
      RECT 187.09 38.41 187.29 65.45 ;
      RECT 185.89 38.41 186.09 65.45 ;
      RECT 184.69 38.41 184.89 65.45 ;
      RECT 183.49 38.41 183.69 65.45 ;
      RECT 182.39 13.78 182.59 24.54 ;
      RECT 182.29 38.41 182.49 65.45 ;
      RECT 181.79 7.04 181.99 9.14 ;
      RECT 181.09 38.41 181.29 65.45 ;
      RECT 180.15 8.84 180.35 9.44 ;
      RECT 179.89 38.41 180.09 65.45 ;
      RECT 179.73 22.31 179.93 24.62 ;
      RECT 179.38 15.39 179.58 16.47 ;
      RECT 179.09 27.45 179.29 37.41 ;
      RECT 177.23 25.27 179.15 25.47 ;
      RECT 177.23 25.67 179.15 25.87 ;
      RECT 178.69 38.41 178.89 65.45 ;
      RECT 177.49 38.41 177.69 65.45 ;
      RECT 177.09 27.45 177.29 37.41 ;
      RECT 176.45 22.31 176.65 24.62 ;
      RECT 176.29 38.41 176.49 65.45 ;
      RECT 175.09 38.41 175.29 65.45 ;
      RECT 173.89 38.41 174.09 65.45 ;
      RECT 173.79 16.5 173.99 24.54 ;
      RECT 172.79 16.5 172.99 24.54 ;
      RECT 172.69 38.41 172.89 65.45 ;
      RECT 171.49 38.41 171.69 65.45 ;
      RECT 170.29 38.41 170.49 65.45 ;
      RECT 170.13 22.31 170.33 24.62 ;
      RECT 169.49 27.45 169.69 37.41 ;
      RECT 167.63 25.27 169.55 25.47 ;
      RECT 167.63 25.67 169.55 25.87 ;
      RECT 169.09 38.41 169.29 65.45 ;
      RECT 167.89 38.41 168.09 65.45 ;
      RECT 167.49 27.45 167.69 37.41 ;
      RECT 167.2 15.39 167.4 16.47 ;
      RECT 166.85 22.31 167.05 24.62 ;
      RECT 166.69 38.41 166.89 65.45 ;
      RECT 166.43 8.84 166.63 9.44 ;
      RECT 165.49 38.41 165.69 65.45 ;
      RECT 164.79 7.04 164.99 9.14 ;
      RECT 164.29 38.41 164.49 65.45 ;
      RECT 164.19 13.78 164.39 24.54 ;
      RECT 163.09 38.41 163.29 65.45 ;
      RECT 161.89 38.41 162.09 65.45 ;
      RECT 160.69 38.41 160.89 65.45 ;
      RECT 159.49 38.41 159.69 65.45 ;
      RECT 158.29 38.41 158.49 65.45 ;
      RECT 157.09 38.41 157.29 65.45 ;
      RECT 155.89 38.41 156.09 65.45 ;
      RECT 154.69 38.41 154.89 65.45 ;
      RECT 152.89 9.34 153.09 22.92 ;
      RECT 149.59 509.8 152.89 510 ;
      RECT 151.99 510.34 152.79 510.94 ;
      RECT 152.09 10.98 152.69 67.63 ;
      RECT 149.61 508.8 152.09 509 ;
      RECT 150.79 510.34 151.59 510.94 ;
      RECT 151.29 22.39 151.49 30.95 ;
      RECT 150.99 31.95 151.39 68.66 ;
      RECT 149.93 510.34 150.39 510.94 ;
      RECT 149.53 52.07 149.73 62.78 ;
      RECT 149.27 7.14 149.47 16.87 ;
      RECT 147.65 16.27 147.85 29.66 ;
      RECT 147.61 52.07 147.81 62.78 ;
      RECT 145.69 52.07 145.89 62.78 ;
      RECT 145.65 23.26 145.85 30.95 ;
      RECT 144.01 7.14 144.21 16.34 ;
      RECT 143.81 16.74 144.01 29.84 ;
      RECT 143.77 52.07 143.97 62.78 ;
      RECT 141.85 52.07 142.05 62.78 ;
      RECT 140.21 24.03 140.41 66.03 ;
      RECT 138.41 12.32 138.61 38.18 ;
      RECT 138.01 7.14 138.21 13.02 ;
      RECT 138.01 16.13 138.21 44.54 ;
      RECT 138.01 44.84 138.21 65.83 ;
      RECT 137.61 13.78 137.81 38.18 ;
      RECT 135.01 13.78 135.21 35.53 ;
      RECT 134.61 7.14 134.81 13.02 ;
      RECT 134.21 12.32 134.41 34.73 ;
      RECT 134.21 35.33 134.41 38.18 ;
      RECT 133.7 32.48 133.9 38.18 ;
      RECT 131.61 35.33 131.81 38.18 ;
      RECT 131.21 7.14 131.41 13.02 ;
      RECT 130.81 13.78 131.01 32.68 ;
      RECT 130.81 34.53 131.01 38.18 ;
      RECT 130.2 34.53 130.4 37.34 ;
      RECT 128.21 13.78 128.41 34.73 ;
      RECT 127.81 7.14 128.01 13.02 ;
      RECT 127.41 12.32 127.61 15.58 ;
      RECT 127.41 35.33 127.61 38.18 ;
      RECT 126.9 32.48 127.1 38.18 ;
      RECT 125.32 34.93 125.52 38.18 ;
      RECT 124.81 35.33 125.01 38.18 ;
      RECT 124.01 15.38 124.21 37.34 ;
      RECT 121.41 510.34 124.21 510.94 ;
      RECT 123.21 67.11 124.01 506.38 ;
      RECT 121.24 67.61 121.71 505.09 ;
      RECT 121.41 13.78 121.61 35.53 ;
      RECT 121.01 7.14 121.21 13.02 ;
      RECT 120.46 67.61 120.94 505.09 ;
      RECT 120.61 12.32 120.81 34.73 ;
      RECT 120.61 35.33 120.81 38.18 ;
      RECT 120.1 32.48 120.3 38.18 ;
      RECT 117.84 67.61 118.31 505.09 ;
      RECT 118.01 35.33 118.21 38.18 ;
      RECT 117.61 7.14 117.81 13.02 ;
      RECT 117.06 67.61 117.54 505.09 ;
      RECT 117.21 13.78 117.41 32.68 ;
      RECT 117.21 34.53 117.41 38.18 ;
      RECT 116.6 34.53 116.8 37.38 ;
      RECT 114.44 67.61 114.91 505.09 ;
      RECT 114.61 13.78 114.81 34.73 ;
      RECT 114.21 7.14 114.41 13.02 ;
      RECT 113.66 67.61 114.14 505.09 ;
      RECT 113.81 12.32 114.01 15.58 ;
      RECT 113.81 35.33 114.01 38.18 ;
      RECT 113.3 32.48 113.5 38.18 ;
      RECT 111.72 34.93 111.92 38.18 ;
      RECT 111.04 67.61 111.51 505.09 ;
      RECT 111.21 35.33 111.41 38.18 ;
      RECT 110.26 67.61 110.74 505.09 ;
      RECT 110.41 15.38 110.61 37.38 ;
      RECT 109.51 509.74 110.61 510.94 ;
      RECT 107.81 509.74 108.91 510.94 ;
      RECT 107.81 13.78 108.01 35.53 ;
      RECT 107.41 7.14 107.61 13.02 ;
      RECT 107.01 12.32 107.21 34.73 ;
      RECT 107.01 35.33 107.21 38.18 ;
      RECT 106.11 509.74 107.21 510.94 ;
      RECT 106.5 32.48 106.7 38.18 ;
      RECT 104.41 509.74 105.51 510.94 ;
      RECT 104.41 35.33 104.61 38.18 ;
      RECT 104.01 7.14 104.21 13.02 ;
      RECT 103.61 13.78 103.81 32.68 ;
      RECT 103.61 34.53 103.81 38.18 ;
      RECT 102.71 509.74 103.81 510.94 ;
      RECT 103 34.53 103.2 37.38 ;
      RECT 101.01 509.74 102.11 510.94 ;
      RECT 101.01 13.78 101.21 34.73 ;
      RECT 100.61 7.14 100.81 13.02 ;
      RECT 100.21 12.32 100.41 15.58 ;
      RECT 100.21 35.33 100.41 38.18 ;
      RECT 99.31 509.74 100.41 510.94 ;
      RECT 99.7 32.48 99.9 38.18 ;
      RECT 97.61 509.74 98.71 510.94 ;
      RECT 98.12 34.93 98.32 38.18 ;
      RECT 97.61 35.33 97.81 38.18 ;
      RECT 96.81 15.38 97.01 37.38 ;
      RECT 95.91 509.74 97.01 510.94 ;
      RECT 94.21 509.74 95.31 510.94 ;
      RECT 94.21 13.78 94.41 38.18 ;
      RECT 93.81 7.14 94.01 13.02 ;
      RECT 93.41 12.32 93.61 38.18 ;
      RECT 92.51 509.74 93.61 510.94 ;
      RECT 92.9 32.51 93.1 38.18 ;
      RECT 90.81 509.74 91.91 510.94 ;
      RECT 90.41 7.14 90.61 13.02 ;
      RECT 90.01 13.78 90.21 32.71 ;
      RECT 89.11 509.74 90.21 510.94 ;
      RECT 0 505.6 88.61 506 ;
      RECT 87.81 510.34 88.61 510.94 ;
      RECT 46.51 507.3 88.1 507.7 ;
      RECT 87.21 6.24 88.01 6.64 ;
      RECT 87.21 10.98 88.01 67.73 ;
      RECT 85.71 38.41 85.91 65.45 ;
      RECT 84.51 38.41 84.71 65.45 ;
      RECT 83.31 38.41 83.51 65.45 ;
      RECT 82.11 38.41 82.31 65.45 ;
      RECT 80.91 38.41 81.11 65.45 ;
      RECT 79.71 38.41 79.91 65.45 ;
      RECT 78.51 38.41 78.71 65.45 ;
      RECT 77.31 38.41 77.51 65.45 ;
      RECT 76.21 13.78 76.41 24.54 ;
      RECT 76.11 38.41 76.31 65.45 ;
      RECT 75.61 7.04 75.81 9.14 ;
      RECT 74.91 38.41 75.11 65.45 ;
      RECT 73.97 8.84 74.17 9.44 ;
      RECT 73.71 38.41 73.91 65.45 ;
      RECT 73.55 22.31 73.75 24.62 ;
      RECT 73.2 15.39 73.4 16.47 ;
      RECT 72.91 27.45 73.11 37.41 ;
      RECT 71.05 25.27 72.97 25.47 ;
      RECT 71.05 25.67 72.97 25.87 ;
      RECT 72.51 38.41 72.71 65.45 ;
      RECT 71.31 38.41 71.51 65.45 ;
      RECT 70.91 27.45 71.11 37.41 ;
      RECT 70.27 22.31 70.47 24.62 ;
      RECT 70.11 38.41 70.31 65.45 ;
      RECT 68.91 38.41 69.11 65.45 ;
      RECT 67.71 38.41 67.91 65.45 ;
      RECT 67.61 16.5 67.81 24.54 ;
      RECT 66.61 16.5 66.81 24.54 ;
      RECT 66.51 38.41 66.71 65.45 ;
      RECT 65.31 38.41 65.51 65.45 ;
      RECT 64.11 38.41 64.31 65.45 ;
      RECT 63.95 22.31 64.15 24.62 ;
      RECT 63.31 27.45 63.51 37.41 ;
      RECT 61.45 25.27 63.37 25.47 ;
      RECT 61.45 25.67 63.37 25.87 ;
      RECT 62.91 38.41 63.11 65.45 ;
      RECT 61.71 38.41 61.91 65.45 ;
      RECT 61.31 27.45 61.51 37.41 ;
      RECT 61.02 15.39 61.22 16.47 ;
      RECT 60.67 22.31 60.87 24.62 ;
      RECT 60.51 38.41 60.71 65.45 ;
      RECT 60.25 8.84 60.45 9.44 ;
      RECT 59.31 38.41 59.51 65.45 ;
      RECT 58.61 7.04 58.81 9.14 ;
      RECT 58.11 38.41 58.31 65.45 ;
      RECT 58.01 13.78 58.21 24.54 ;
      RECT 56.91 38.41 57.11 65.45 ;
      RECT 55.71 38.41 55.91 65.45 ;
      RECT 54.51 38.41 54.71 65.45 ;
      RECT 53.31 38.41 53.51 65.45 ;
      RECT 52.11 38.41 52.31 65.45 ;
      RECT 50.91 38.41 51.11 65.45 ;
      RECT 49.71 38.41 49.91 65.45 ;
      RECT 48.51 38.41 48.71 65.45 ;
      RECT 47.31 57.02 47.51 63.45 ;
      RECT 46.11 38.41 46.31 65.45 ;
      RECT 44.91 38.41 45.11 65.45 ;
      RECT 43.71 38.41 43.91 65.45 ;
      RECT 42.51 38.41 42.71 65.45 ;
      RECT 41.31 38.41 41.51 65.45 ;
      RECT 40.11 38.41 40.31 65.45 ;
      RECT 38.91 38.41 39.11 65.45 ;
      RECT 37.71 38.41 37.91 65.45 ;
      RECT 36.61 13.78 36.81 24.54 ;
      RECT 36.51 38.41 36.71 65.45 ;
      RECT 36.01 7.04 36.21 9.14 ;
      RECT 35.31 38.41 35.51 65.45 ;
      RECT 34.37 8.84 34.57 9.44 ;
      RECT 34.11 38.41 34.31 65.45 ;
      RECT 33.95 22.31 34.15 24.62 ;
      RECT 33.6 15.39 33.8 16.47 ;
      RECT 33.31 27.45 33.51 37.41 ;
      RECT 31.45 25.27 33.37 25.47 ;
      RECT 31.45 25.67 33.37 25.87 ;
      RECT 32.91 38.41 33.11 65.45 ;
      RECT 31.71 38.41 31.91 65.45 ;
      RECT 31.31 27.45 31.51 37.41 ;
      RECT 30.67 22.31 30.87 24.62 ;
      RECT 30.51 38.41 30.71 65.45 ;
      RECT 29.31 38.41 29.51 65.45 ;
      RECT 28.11 38.41 28.31 65.45 ;
      RECT 28.01 16.5 28.21 24.54 ;
      RECT 27.01 16.5 27.21 24.54 ;
      RECT 26.91 38.41 27.11 65.45 ;
      RECT 25.71 38.41 25.91 65.45 ;
      RECT 24.51 38.41 24.71 65.45 ;
      RECT 24.35 22.31 24.55 24.62 ;
      RECT 23.71 27.45 23.91 37.41 ;
      RECT 21.85 25.27 23.77 25.47 ;
      RECT 21.85 25.67 23.77 25.87 ;
      RECT 23.31 38.41 23.51 65.45 ;
      RECT 22.11 38.41 22.31 65.45 ;
      RECT 21.71 27.45 21.91 37.41 ;
      RECT 21.42 15.39 21.62 16.47 ;
      RECT 21.07 22.31 21.27 24.62 ;
      RECT 20.91 38.41 21.11 65.45 ;
      RECT 20.65 8.84 20.85 9.44 ;
      RECT 19.71 38.41 19.91 65.45 ;
      RECT 18.51 38.41 18.71 65.45 ;
      RECT 18.41 13.78 18.61 24.54 ;
      RECT 17.31 38.41 17.51 65.45 ;
      RECT 16.11 38.41 16.31 65.45 ;
      RECT 14.91 38.41 15.11 65.45 ;
      RECT 13.71 38.41 13.91 65.45 ;
      RECT 12.51 38.41 12.71 65.45 ;
      RECT 11.31 38.41 11.51 65.45 ;
      RECT 10.11 38.41 10.31 65.45 ;
      RECT 8.91 38.41 9.11 65.45 ;
      RECT 0 7.94 6.84 9.14 ;
      RECT 0 17.26 6.84 18.46 ;
      RECT 0 25.81 6.84 27.81 ;
      RECT 0 35.91 6.84 36.91 ;
      RECT 0 50.24 6.84 51.24 ;
      RECT 0 57.02 6.84 58.02 ;
      RECT 0 60.6 6.84 61.6 ;
      RECT 0 62.45 6.84 63.45 ;
    LAYER M4 ;
      RECT 232.39 3.12 233.19 514.06 ;
      RECT 231.19 3.12 231.99 514.06 ;
      RECT 231.19 510.34 233.39 510.74 ;
      RECT 232.39 506.6 234.36 508.6 ;
      RECT 232.39 502.66 234.36 503.46 ;
      RECT 232.39 499.26 234.36 500.06 ;
      RECT 232.39 495.86 234.36 496.66 ;
      RECT 232.39 492.46 234.36 493.26 ;
      RECT 232.39 489.06 234.36 489.86 ;
      RECT 232.39 485.66 234.36 486.46 ;
      RECT 232.39 482.26 234.36 483.06 ;
      RECT 232.39 478.86 234.36 479.66 ;
      RECT 232.39 475.46 234.36 476.26 ;
      RECT 232.39 472.06 234.36 472.86 ;
      RECT 232.39 468.66 234.36 469.46 ;
      RECT 232.39 465.26 234.36 466.06 ;
      RECT 232.39 461.86 234.36 462.66 ;
      RECT 232.39 458.46 234.36 459.26 ;
      RECT 232.39 455.06 234.36 455.86 ;
      RECT 232.39 451.66 234.36 452.46 ;
      RECT 232.39 448.26 234.36 449.06 ;
      RECT 232.39 444.86 234.36 445.66 ;
      RECT 232.39 441.46 234.36 442.26 ;
      RECT 232.39 438.06 234.36 438.86 ;
      RECT 232.39 434.66 234.36 435.46 ;
      RECT 232.39 431.26 234.36 432.06 ;
      RECT 232.39 427.86 234.36 428.66 ;
      RECT 232.39 424.46 234.36 425.26 ;
      RECT 232.39 421.06 234.36 421.86 ;
      RECT 232.39 417.66 234.36 418.46 ;
      RECT 232.39 414.26 234.36 415.06 ;
      RECT 232.39 410.86 234.36 411.66 ;
      RECT 232.39 407.46 234.36 408.26 ;
      RECT 232.39 404.06 234.36 404.86 ;
      RECT 232.39 400.66 234.36 401.46 ;
      RECT 232.39 397.26 234.36 398.06 ;
      RECT 232.39 393.86 234.36 394.66 ;
      RECT 232.39 390.46 234.36 391.26 ;
      RECT 232.39 387.06 234.36 387.86 ;
      RECT 232.39 383.66 234.36 384.46 ;
      RECT 232.39 380.26 234.36 381.06 ;
      RECT 232.39 376.86 234.36 377.66 ;
      RECT 232.39 373.46 234.36 374.26 ;
      RECT 232.39 370.06 234.36 370.86 ;
      RECT 232.39 366.66 234.36 367.46 ;
      RECT 232.39 363.26 234.36 364.06 ;
      RECT 232.39 359.86 234.36 360.66 ;
      RECT 232.39 356.46 234.36 357.26 ;
      RECT 232.39 353.06 234.36 353.86 ;
      RECT 232.39 349.66 234.36 350.46 ;
      RECT 232.39 346.26 234.36 347.06 ;
      RECT 232.39 342.86 234.36 343.66 ;
      RECT 232.39 339.46 234.36 340.26 ;
      RECT 232.39 336.06 234.36 336.86 ;
      RECT 232.39 332.66 234.36 333.46 ;
      RECT 232.39 329.26 234.36 330.06 ;
      RECT 232.39 325.86 234.36 326.66 ;
      RECT 232.39 322.46 234.36 323.26 ;
      RECT 232.39 319.06 234.36 319.86 ;
      RECT 232.39 315.66 234.36 316.46 ;
      RECT 232.39 312.26 234.36 313.06 ;
      RECT 232.39 308.86 234.36 309.66 ;
      RECT 232.39 305.46 234.36 306.26 ;
      RECT 232.39 302.06 234.36 302.86 ;
      RECT 232.39 298.66 234.36 299.46 ;
      RECT 232.39 295.26 234.36 296.06 ;
      RECT 232.39 291.86 234.36 292.66 ;
      RECT 232.39 288.46 234.36 289.26 ;
      RECT 232.39 285.06 234.36 285.86 ;
      RECT 232.39 281.66 234.36 282.46 ;
      RECT 232.39 278.26 234.36 279.06 ;
      RECT 232.39 274.86 234.36 275.66 ;
      RECT 232.39 271.46 234.36 272.26 ;
      RECT 232.39 268.06 234.36 268.86 ;
      RECT 232.39 264.66 234.36 265.46 ;
      RECT 232.39 261.26 234.36 262.06 ;
      RECT 232.39 257.86 234.36 258.66 ;
      RECT 232.39 254.46 234.36 255.26 ;
      RECT 232.39 251.06 234.36 251.86 ;
      RECT 232.39 247.66 234.36 248.46 ;
      RECT 232.39 244.26 234.36 245.06 ;
      RECT 232.39 240.86 234.36 241.66 ;
      RECT 232.39 237.46 234.36 238.26 ;
      RECT 232.39 234.06 234.36 234.86 ;
      RECT 232.39 230.66 234.36 231.46 ;
      RECT 232.39 227.26 234.36 228.06 ;
      RECT 232.39 223.86 234.36 224.66 ;
      RECT 232.39 220.46 234.36 221.26 ;
      RECT 232.39 217.06 234.36 217.86 ;
      RECT 232.39 213.66 234.36 214.46 ;
      RECT 232.39 210.26 234.36 211.06 ;
      RECT 232.39 206.86 234.36 207.66 ;
      RECT 232.39 203.46 234.36 204.26 ;
      RECT 232.39 200.06 234.36 200.86 ;
      RECT 232.39 196.66 234.36 197.46 ;
      RECT 232.39 193.26 234.36 194.06 ;
      RECT 232.39 189.86 234.36 190.66 ;
      RECT 232.39 186.46 234.36 187.26 ;
      RECT 232.39 183.06 234.36 183.86 ;
      RECT 232.39 179.66 234.36 180.46 ;
      RECT 232.39 176.26 234.36 177.06 ;
      RECT 232.39 172.86 234.36 173.66 ;
      RECT 232.39 169.46 234.36 170.26 ;
      RECT 232.39 166.06 234.36 166.86 ;
      RECT 232.39 162.66 234.36 163.46 ;
      RECT 232.39 159.26 234.36 160.06 ;
      RECT 232.39 155.86 234.36 156.66 ;
      RECT 232.39 152.46 234.36 153.26 ;
      RECT 232.39 149.06 234.36 149.86 ;
      RECT 232.39 145.66 234.36 146.46 ;
      RECT 232.39 142.26 234.36 143.06 ;
      RECT 232.39 138.86 234.36 139.66 ;
      RECT 232.39 135.46 234.36 136.26 ;
      RECT 232.39 132.06 234.36 132.86 ;
      RECT 232.39 128.66 234.36 129.46 ;
      RECT 232.39 125.26 234.36 126.06 ;
      RECT 232.39 121.86 234.36 122.66 ;
      RECT 232.39 118.46 234.36 119.26 ;
      RECT 232.39 115.06 234.36 115.86 ;
      RECT 232.39 111.66 234.36 112.46 ;
      RECT 232.39 108.26 234.36 109.06 ;
      RECT 232.39 104.86 234.36 105.66 ;
      RECT 232.39 101.46 234.36 102.26 ;
      RECT 232.39 98.06 234.36 98.86 ;
      RECT 232.39 94.66 234.36 95.46 ;
      RECT 232.39 91.26 234.36 92.06 ;
      RECT 232.39 87.86 234.36 88.66 ;
      RECT 232.39 84.46 234.36 85.26 ;
      RECT 232.39 81.06 234.36 81.86 ;
      RECT 232.39 77.66 234.36 78.46 ;
      RECT 232.39 74.26 234.36 75.06 ;
      RECT 232.39 70.86 234.36 71.66 ;
      RECT 231.19 3.12 233.19 67.05 ;
      RECT 231.19 54.22 234.36 55.22 ;
      RECT 231.19 41.29 234.36 42.29 ;
      RECT 231.19 39.44 234.36 40.44 ;
      RECT 231.19 32.98 234.36 33.98 ;
      RECT 231.19 31.13 234.36 32.13 ;
      RECT 231.19 21.41 234.36 22.21 ;
      RECT 231.19 12.64 234.36 13.74 ;
      RECT 233.76 505.6 234.36 506 ;
      RECT 233.76 504.36 234.16 506 ;
      RECT 233.76 504.36 234.36 505.16 ;
      RECT 228.79 510.34 230.79 517.18 ;
      RECT 229.99 0 230.79 517.18 ;
      RECT 228.79 7.44 229.59 517.18 ;
      RECT 228.81 0 230.79 67.05 ;
      RECT 227.59 3.12 228.39 514.06 ;
      RECT 226.39 7.44 227.19 514.06 ;
      RECT 226.39 510.34 228.39 510.74 ;
      RECT 226.41 3.12 228.39 67.05 ;
      RECT 223.99 510.34 225.99 517.18 ;
      RECT 225.19 0 225.99 517.18 ;
      RECT 223.99 7.44 224.79 517.18 ;
      RECT 224.01 0 225.99 67.05 ;
      RECT 222.79 3.12 223.59 514.06 ;
      RECT 221.59 3.12 222.39 514.06 ;
      RECT 221.59 510.34 223.59 510.74 ;
      RECT 221.59 3.12 223.59 67.05 ;
      RECT 219.19 510.34 221.19 517.18 ;
      RECT 220.39 0 221.19 517.18 ;
      RECT 219.19 7.44 219.99 517.18 ;
      RECT 219.21 0 221.19 67.05 ;
      RECT 217.99 3.12 218.79 514.06 ;
      RECT 216.79 7.44 217.59 514.06 ;
      RECT 216.79 510.34 218.79 510.74 ;
      RECT 217.29 3.12 218.79 67.05 ;
      RECT 214.39 510.34 216.39 517.18 ;
      RECT 215.59 7.44 216.39 517.18 ;
      RECT 214.39 7.44 215.19 517.18 ;
      RECT 214.89 0 215.89 67.05 ;
      RECT 213.19 7.44 213.99 514.06 ;
      RECT 211.99 7.44 212.79 514.06 ;
      RECT 211.99 510.34 213.99 510.74 ;
      RECT 212.59 3.12 213.39 67.05 ;
      RECT 209.59 510.34 211.59 517.18 ;
      RECT 210.79 7.44 211.59 517.18 ;
      RECT 209.59 7.44 210.39 517.18 ;
      RECT 210.09 0 211.09 67.05 ;
      RECT 208.39 7.44 209.19 514.06 ;
      RECT 207.19 3.12 207.99 514.06 ;
      RECT 207.19 510.34 209.19 510.74 ;
      RECT 207.19 3.12 208.69 67.05 ;
      RECT 204.79 510.34 206.79 517.18 ;
      RECT 205.99 7.44 206.79 517.18 ;
      RECT 204.79 0 205.59 517.18 ;
      RECT 204.79 0 206.76 67.05 ;
      RECT 203.59 3.12 204.39 514.06 ;
      RECT 202.39 3.12 203.19 514.06 ;
      RECT 202.39 510.34 204.39 510.74 ;
      RECT 202.39 3.12 204.39 67.05 ;
      RECT 199.99 510.34 201.99 517.18 ;
      RECT 201.19 7.44 201.99 517.18 ;
      RECT 199.99 0 200.79 517.18 ;
      RECT 199.99 0 201.97 67.05 ;
      RECT 198.79 7.44 199.59 514.06 ;
      RECT 197.59 3.12 198.39 514.06 ;
      RECT 197.59 510.34 199.59 510.74 ;
      RECT 197.59 3.12 199.57 67.05 ;
      RECT 195.19 510.34 197.19 517.18 ;
      RECT 196.39 7.44 197.19 517.18 ;
      RECT 195.19 0 195.99 517.18 ;
      RECT 195.19 0 197.17 67.05 ;
      RECT 193.99 3.12 194.79 514.06 ;
      RECT 192.79 65.72 193.59 514.06 ;
      RECT 191.59 3.12 192.39 514.06 ;
      RECT 191.59 510.34 194.79 510.74 ;
      RECT 193.39 3.12 194.79 67.05 ;
      RECT 191.59 3.12 192.99 67.05 ;
      RECT 189.19 510.34 191.19 517.18 ;
      RECT 190.39 0 191.19 517.18 ;
      RECT 189.19 7.44 189.99 517.18 ;
      RECT 189.21 0 191.19 67.05 ;
      RECT 187.99 3.12 188.79 514.06 ;
      RECT 186.79 7.44 187.59 514.06 ;
      RECT 186.79 510.34 188.79 510.74 ;
      RECT 186.81 3.12 188.79 67.05 ;
      RECT 184.39 510.34 186.39 517.18 ;
      RECT 185.59 0 186.39 517.18 ;
      RECT 184.39 7.44 185.19 517.18 ;
      RECT 184.41 0 186.39 67.05 ;
      RECT 183.19 3.12 183.99 514.06 ;
      RECT 181.99 3.12 182.79 514.06 ;
      RECT 181.99 510.34 183.99 510.74 ;
      RECT 181.99 3.12 183.99 67.05 ;
      RECT 179.59 510.34 181.59 517.18 ;
      RECT 180.79 0 181.59 517.18 ;
      RECT 179.59 7.44 180.39 517.18 ;
      RECT 179.62 0 181.59 67.05 ;
      RECT 178.39 3.12 179.19 514.06 ;
      RECT 177.19 7.44 177.99 514.06 ;
      RECT 177.19 510.34 179.19 510.74 ;
      RECT 177.69 3.12 179.19 67.05 ;
      RECT 174.79 510.34 176.79 517.18 ;
      RECT 175.99 7.44 176.79 517.18 ;
      RECT 174.79 7.44 175.59 517.18 ;
      RECT 175.29 0 176.29 67.05 ;
      RECT 173.59 7.44 174.39 514.06 ;
      RECT 172.39 7.44 173.19 514.06 ;
      RECT 172.39 510.34 174.39 510.74 ;
      RECT 172.99 3.12 173.79 67.05 ;
      RECT 169.99 510.34 171.99 517.18 ;
      RECT 171.19 7.44 171.99 517.18 ;
      RECT 169.99 7.44 170.79 517.18 ;
      RECT 170.49 0 171.49 67.05 ;
      RECT 168.79 7.44 169.59 514.06 ;
      RECT 167.59 3.12 168.39 514.06 ;
      RECT 167.59 510.34 169.59 510.74 ;
      RECT 167.59 3.12 169.09 67.05 ;
      RECT 165.19 510.34 167.19 517.18 ;
      RECT 166.39 7.44 167.19 517.18 ;
      RECT 165.19 0 165.99 517.18 ;
      RECT 165.19 0 167.16 67.05 ;
      RECT 163.99 3.12 164.79 514.06 ;
      RECT 162.79 3.12 163.59 514.06 ;
      RECT 162.79 510.34 164.79 510.74 ;
      RECT 162.79 3.12 164.79 67.05 ;
      RECT 160.39 510.34 162.39 517.18 ;
      RECT 161.59 7.44 162.39 517.18 ;
      RECT 160.39 0 161.19 517.18 ;
      RECT 160.39 0 162.37 67.05 ;
      RECT 159.19 7.44 159.99 514.06 ;
      RECT 157.99 3.12 158.79 514.06 ;
      RECT 157.99 510.34 159.99 510.74 ;
      RECT 157.99 3.12 159.97 67.05 ;
      RECT 155.59 510.34 157.59 517.18 ;
      RECT 156.79 7.44 157.59 517.18 ;
      RECT 155.59 0 156.39 517.18 ;
      RECT 155.59 0 157.57 67.05 ;
      RECT 154.39 3.12 155.19 514.06 ;
      RECT 153.19 8.19 153.99 514.06 ;
      RECT 153.19 510.34 155.19 510.74 ;
      RECT 153.89 3.12 155.19 67.05 ;
      RECT 150.79 8.19 151.59 514.06 ;
      RECT 149.93 8.19 150.39 514.06 ;
      RECT 150.29 3.12 150.89 67.13 ;
      RECT 148.01 8.19 149.33 517.18 ;
      RECT 148.01 0 148.87 517.18 ;
      RECT 144.17 8.19 145.49 517.18 ;
      RECT 145.01 0 145.61 8.59 ;
      RECT 142.25 8.19 143.57 514.06 ;
      RECT 142.62 3.12 143.57 514.06 ;
      RECT 138.41 8.19 141.65 517.18 ;
      RECT 138.83 0 140.83 517.18 ;
      RECT 135.01 67.73 137.81 514.06 ;
      RECT 136.71 8.19 137.81 514.06 ;
      RECT 133.31 67.73 137.81 68.83 ;
      RECT 133.31 66.63 134.41 68.83 ;
      RECT 135.01 8.19 137.81 64.43 ;
      RECT 135.43 3.12 137.39 64.43 ;
      RECT 131.61 69.43 134.41 517.18 ;
      RECT 131.61 8.19 132.71 517.18 ;
      RECT 135.01 65.03 136.11 67.13 ;
      RECT 131.61 65.03 136.11 66.03 ;
      RECT 131.61 8.19 134.41 66.03 ;
      RECT 132.03 0 133.99 66.03 ;
      RECT 128.21 67.73 131.01 514.06 ;
      RECT 129.91 8.19 131.01 514.06 ;
      RECT 126.51 67.73 131.01 68.83 ;
      RECT 126.51 66.63 127.61 68.83 ;
      RECT 128.21 8.19 131.01 64.43 ;
      RECT 128.63 3.12 130.59 64.43 ;
      RECT 124.81 69.43 127.61 517.18 ;
      RECT 124.81 8.19 125.91 517.18 ;
      RECT 128.21 65.03 129.31 67.13 ;
      RECT 124.81 65.03 129.31 66.03 ;
      RECT 124.81 8.19 127.61 66.03 ;
      RECT 125.21 0 127.19 66.03 ;
      RECT 121.41 67.73 124.21 514.06 ;
      RECT 123.11 8.19 124.21 514.06 ;
      RECT 119.71 67.73 124.21 68.83 ;
      RECT 119.71 66.63 120.81 68.83 ;
      RECT 121.41 8.19 124.21 64.43 ;
      RECT 121.83 3.12 123.81 64.43 ;
      RECT 118.01 69.43 120.81 517.18 ;
      RECT 118.01 8.19 119.11 517.18 ;
      RECT 121.41 65.03 122.51 67.13 ;
      RECT 118.01 65.03 122.51 66.03 ;
      RECT 118.01 8.19 120.81 66.03 ;
      RECT 118.43 0 120.39 66.03 ;
      RECT 114.61 67.73 117.41 514.06 ;
      RECT 116.31 8.19 117.41 514.06 ;
      RECT 112.91 67.73 117.41 68.83 ;
      RECT 112.91 66.63 114.01 68.83 ;
      RECT 114.61 8.19 117.41 64.43 ;
      RECT 115.03 3.12 116.99 64.43 ;
      RECT 111.21 69.43 114.01 517.18 ;
      RECT 111.21 8.19 112.31 517.18 ;
      RECT 114.61 65.03 115.71 67.13 ;
      RECT 111.21 65.03 115.71 66.03 ;
      RECT 111.21 8.19 114.01 66.03 ;
      RECT 111.61 0 113.59 66.03 ;
      RECT 109.51 8.19 110.61 514.06 ;
      RECT 107.81 8.19 110.61 64.43 ;
      RECT 108.23 3.12 110.21 64.43 ;
      RECT 107.81 65.03 108.91 517.18 ;
      RECT 104.41 8.19 105.51 517.18 ;
      RECT 104.41 65.03 108.91 66.03 ;
      RECT 104.41 8.19 107.21 66.03 ;
      RECT 104.83 0 106.79 66.03 ;
      RECT 102.71 8.19 103.81 514.06 ;
      RECT 101.01 8.19 103.81 64.43 ;
      RECT 101.43 3.12 103.39 64.43 ;
      RECT 101.01 65.03 102.11 517.18 ;
      RECT 97.61 8.19 98.71 517.18 ;
      RECT 97.61 65.03 102.11 66.03 ;
      RECT 97.61 8.19 100.41 66.03 ;
      RECT 98.01 0 99.99 66.03 ;
      RECT 95.91 8.19 97.01 514.06 ;
      RECT 94.21 8.19 97.01 64.43 ;
      RECT 94.63 3.12 96.61 64.43 ;
      RECT 94.21 65.03 95.31 517.18 ;
      RECT 90.81 8.19 91.91 517.18 ;
      RECT 90.81 65.03 95.31 66.03 ;
      RECT 90.81 8.19 93.61 66.03 ;
      RECT 91.23 0 93.19 66.03 ;
      RECT 89.11 8.19 90.21 514.06 ;
      RECT 88.81 3.12 89.79 64.43 ;
      RECT 88.61 6.24 89.79 64.43 ;
      RECT 87.81 67.13 88.61 517.18 ;
      RECT 87.21 0 88.01 68.47 ;
      RECT 86.61 68.94 87.41 514.06 ;
      RECT 85.41 3.12 86.21 514.06 ;
      RECT 85.41 510.34 87.41 510.74 ;
      RECT 85.41 3.12 86.61 67.05 ;
      RECT 85.41 3.12 86.71 7.44 ;
      RECT 83.01 510.34 85.01 517.18 ;
      RECT 84.21 0 85.01 517.18 ;
      RECT 83.01 7.44 83.81 517.18 ;
      RECT 83.03 0 85.01 67.05 ;
      RECT 81.81 3.12 82.61 514.06 ;
      RECT 80.61 7.44 81.41 514.06 ;
      RECT 80.61 510.34 82.61 510.74 ;
      RECT 80.63 3.12 82.61 67.05 ;
      RECT 78.21 510.34 80.21 517.18 ;
      RECT 79.41 0 80.21 517.18 ;
      RECT 78.21 7.44 79.01 517.18 ;
      RECT 78.23 0 80.21 67.05 ;
      RECT 77.01 3.12 77.81 514.06 ;
      RECT 75.81 3.12 76.61 514.06 ;
      RECT 75.81 510.34 77.81 510.74 ;
      RECT 75.81 3.12 77.81 67.05 ;
      RECT 73.41 510.34 75.41 517.18 ;
      RECT 74.61 0 75.41 517.18 ;
      RECT 73.41 7.44 74.21 517.18 ;
      RECT 73.44 0 75.41 67.05 ;
      RECT 72.21 3.12 73.01 514.06 ;
      RECT 71.01 7.44 71.81 514.06 ;
      RECT 71.01 510.34 73.01 510.74 ;
      RECT 71.51 3.12 73.01 67.05 ;
      RECT 68.61 510.34 70.61 517.18 ;
      RECT 69.81 7.44 70.61 517.18 ;
      RECT 68.61 7.44 69.41 517.18 ;
      RECT 69.11 0 70.11 67.05 ;
      RECT 67.41 7.44 68.21 514.06 ;
      RECT 66.21 7.44 67.01 514.06 ;
      RECT 66.21 510.34 68.21 510.74 ;
      RECT 66.81 3.12 67.61 67.05 ;
      RECT 63.81 510.34 65.81 517.18 ;
      RECT 65.01 7.44 65.81 517.18 ;
      RECT 63.81 7.44 64.61 517.18 ;
      RECT 64.31 0 65.31 67.05 ;
      RECT 62.61 7.44 63.41 514.06 ;
      RECT 61.41 3.12 62.21 514.06 ;
      RECT 61.41 510.34 63.41 510.74 ;
      RECT 61.41 3.12 62.91 67.05 ;
      RECT 59.01 510.34 61.01 517.18 ;
      RECT 60.21 7.44 61.01 517.18 ;
      RECT 59.01 0 59.81 517.18 ;
      RECT 59.01 0 60.98 67.05 ;
      RECT 57.81 3.12 58.61 514.06 ;
      RECT 56.61 3.12 57.41 514.06 ;
      RECT 56.61 510.34 58.61 510.74 ;
      RECT 56.61 3.12 58.61 67.05 ;
      RECT 54.21 510.34 56.21 517.18 ;
      RECT 55.41 7.44 56.21 517.18 ;
      RECT 54.21 0 55.01 517.18 ;
      RECT 54.21 0 56.19 67.05 ;
      RECT 53.01 7.44 53.81 514.06 ;
      RECT 51.81 3.12 52.61 514.06 ;
      RECT 51.81 510.34 53.81 510.74 ;
      RECT 51.81 3.12 53.79 67.05 ;
      RECT 49.41 510.34 51.41 517.18 ;
      RECT 50.61 7.44 51.41 517.18 ;
      RECT 49.41 0 50.21 517.18 ;
      RECT 49.41 0 51.39 67.05 ;
      RECT 48.21 3.12 49.01 514.06 ;
      RECT 47.01 65.72 47.81 514.06 ;
      RECT 45.81 3.12 46.61 514.06 ;
      RECT 45.81 510.34 49.01 510.74 ;
      RECT 47.61 3.12 49.01 67.05 ;
      RECT 45.81 3.12 47.21 67.05 ;
      RECT 43.41 510.34 45.41 517.18 ;
      RECT 44.61 0 45.41 517.18 ;
      RECT 43.41 7.44 44.21 517.18 ;
      RECT 43.43 0 45.41 67.05 ;
      RECT 42.21 3.12 43.01 514.06 ;
      RECT 41.01 7.44 41.81 514.06 ;
      RECT 41.01 510.34 43.01 510.74 ;
      RECT 41.03 3.12 43.01 67.05 ;
      RECT 38.61 510.34 40.61 517.18 ;
      RECT 39.81 0 40.61 517.18 ;
      RECT 38.61 7.44 39.41 517.18 ;
      RECT 38.63 0 40.61 67.05 ;
      RECT 37.41 3.12 38.21 514.06 ;
      RECT 36.21 3.12 37.01 514.06 ;
      RECT 36.21 510.34 38.21 510.74 ;
      RECT 36.21 3.12 38.21 67.05 ;
      RECT 33.81 510.34 35.81 517.18 ;
      RECT 35.01 0 35.81 517.18 ;
      RECT 33.81 7.44 34.61 517.18 ;
      RECT 33.84 0 35.81 67.05 ;
      RECT 32.61 3.12 33.41 514.06 ;
      RECT 31.41 7.44 32.21 514.06 ;
      RECT 31.41 510.34 33.41 510.74 ;
      RECT 31.91 3.12 33.41 67.05 ;
      RECT 29.01 510.34 31.01 517.18 ;
      RECT 30.21 7.44 31.01 517.18 ;
      RECT 29.01 7.44 29.81 517.18 ;
      RECT 29.51 0 30.51 67.05 ;
      RECT 27.81 7.44 28.61 514.06 ;
      RECT 26.61 7.44 27.41 514.06 ;
      RECT 26.61 510.34 28.61 510.74 ;
      RECT 27.21 3.12 28.01 67.05 ;
      RECT 24.21 510.34 26.21 517.18 ;
      RECT 25.41 7.44 26.21 517.18 ;
      RECT 24.21 7.44 25.01 517.18 ;
      RECT 24.71 0 25.71 67.05 ;
      RECT 23.01 7.44 23.81 514.06 ;
      RECT 21.81 3.12 22.61 514.06 ;
      RECT 21.81 510.34 23.81 510.74 ;
      RECT 21.81 3.12 23.31 67.05 ;
      RECT 19.41 510.34 21.41 517.18 ;
      RECT 20.61 0 21.41 517.18 ;
      RECT 19.41 7.44 20.21 517.18 ;
      RECT 19.81 0 21.41 67.05 ;
      RECT 18.21 7.44 19.01 514.06 ;
      RECT 17.01 3.12 17.81 514.06 ;
      RECT 17.01 510.34 19.01 510.74 ;
      RECT 17.01 3.12 18.41 67.05 ;
      RECT 14.61 510.34 16.61 517.18 ;
      RECT 15.81 7.44 16.61 517.18 ;
      RECT 14.61 0 15.41 517.18 ;
      RECT 14.61 0 16.59 67.05 ;
      RECT 13.41 7.44 14.21 514.06 ;
      RECT 12.21 3.12 13.01 514.06 ;
      RECT 12.21 510.34 14.21 510.74 ;
      RECT 12.21 3.12 14.19 67.05 ;
      RECT 9.81 510.34 11.81 517.18 ;
      RECT 11.01 7.44 11.81 517.18 ;
      RECT 9.81 0 10.61 517.18 ;
      RECT 9.81 0 11.79 67.05 ;
      RECT 8.61 3.12 9.41 514.06 ;
      RECT 7.41 3.12 8.21 514.06 ;
      RECT 7.21 510.34 9.41 510.74 ;
      RECT 6.24 506.6 8.21 508.6 ;
      RECT 6.24 502.66 8.21 503.46 ;
      RECT 6.24 499.26 8.21 500.06 ;
      RECT 6.24 495.86 8.21 496.66 ;
      RECT 6.24 492.46 8.21 493.26 ;
      RECT 6.24 489.06 8.21 489.86 ;
      RECT 6.24 485.66 8.21 486.46 ;
      RECT 6.24 482.26 8.21 483.06 ;
      RECT 6.24 478.86 8.21 479.66 ;
      RECT 6.24 475.46 8.21 476.26 ;
      RECT 6.24 472.06 8.21 472.86 ;
      RECT 6.24 468.66 8.21 469.46 ;
      RECT 6.24 465.26 8.21 466.06 ;
      RECT 6.24 461.86 8.21 462.66 ;
      RECT 6.24 458.46 8.21 459.26 ;
      RECT 6.24 455.06 8.21 455.86 ;
      RECT 6.24 451.66 8.21 452.46 ;
      RECT 6.24 448.26 8.21 449.06 ;
      RECT 6.24 444.86 8.21 445.66 ;
      RECT 6.24 441.46 8.21 442.26 ;
      RECT 6.24 438.06 8.21 438.86 ;
      RECT 6.24 434.66 8.21 435.46 ;
      RECT 6.24 431.26 8.21 432.06 ;
      RECT 6.24 427.86 8.21 428.66 ;
      RECT 6.24 424.46 8.21 425.26 ;
      RECT 6.24 421.06 8.21 421.86 ;
      RECT 6.24 417.66 8.21 418.46 ;
      RECT 6.24 414.26 8.21 415.06 ;
      RECT 6.24 410.86 8.21 411.66 ;
      RECT 6.24 407.46 8.21 408.26 ;
      RECT 6.24 404.06 8.21 404.86 ;
      RECT 6.24 400.66 8.21 401.46 ;
      RECT 6.24 397.26 8.21 398.06 ;
      RECT 6.24 393.86 8.21 394.66 ;
      RECT 6.24 390.46 8.21 391.26 ;
      RECT 6.24 387.06 8.21 387.86 ;
      RECT 6.24 383.66 8.21 384.46 ;
      RECT 6.24 380.26 8.21 381.06 ;
      RECT 6.24 376.86 8.21 377.66 ;
      RECT 6.24 373.46 8.21 374.26 ;
      RECT 6.24 370.06 8.21 370.86 ;
      RECT 6.24 366.66 8.21 367.46 ;
      RECT 6.24 363.26 8.21 364.06 ;
      RECT 6.24 359.86 8.21 360.66 ;
      RECT 6.24 356.46 8.21 357.26 ;
      RECT 6.24 353.06 8.21 353.86 ;
      RECT 6.24 349.66 8.21 350.46 ;
      RECT 6.24 346.26 8.21 347.06 ;
      RECT 6.24 342.86 8.21 343.66 ;
      RECT 6.24 339.46 8.21 340.26 ;
      RECT 6.24 336.06 8.21 336.86 ;
      RECT 6.24 332.66 8.21 333.46 ;
      RECT 6.24 329.26 8.21 330.06 ;
      RECT 6.24 325.86 8.21 326.66 ;
      RECT 6.24 322.46 8.21 323.26 ;
      RECT 6.24 319.06 8.21 319.86 ;
      RECT 6.24 315.66 8.21 316.46 ;
      RECT 6.24 312.26 8.21 313.06 ;
      RECT 6.24 308.86 8.21 309.66 ;
      RECT 6.24 305.46 8.21 306.26 ;
      RECT 6.24 302.06 8.21 302.86 ;
      RECT 6.24 298.66 8.21 299.46 ;
      RECT 6.24 295.26 8.21 296.06 ;
      RECT 6.24 291.86 8.21 292.66 ;
      RECT 6.24 288.46 8.21 289.26 ;
      RECT 6.24 285.06 8.21 285.86 ;
      RECT 6.24 281.66 8.21 282.46 ;
      RECT 6.24 278.26 8.21 279.06 ;
      RECT 6.24 274.86 8.21 275.66 ;
      RECT 6.24 271.46 8.21 272.26 ;
      RECT 6.24 268.06 8.21 268.86 ;
      RECT 6.24 264.66 8.21 265.46 ;
      RECT 6.24 261.26 8.21 262.06 ;
      RECT 6.24 257.86 8.21 258.66 ;
      RECT 6.24 254.46 8.21 255.26 ;
      RECT 6.24 251.06 8.21 251.86 ;
      RECT 6.24 247.66 8.21 248.46 ;
      RECT 6.24 244.26 8.21 245.06 ;
      RECT 6.24 240.86 8.21 241.66 ;
      RECT 6.24 237.46 8.21 238.26 ;
      RECT 6.24 234.06 8.21 234.86 ;
      RECT 6.24 230.66 8.21 231.46 ;
      RECT 6.24 227.26 8.21 228.06 ;
      RECT 6.24 223.86 8.21 224.66 ;
      RECT 6.24 220.46 8.21 221.26 ;
      RECT 6.24 217.06 8.21 217.86 ;
      RECT 6.24 213.66 8.21 214.46 ;
      RECT 6.24 210.26 8.21 211.06 ;
      RECT 6.24 206.86 8.21 207.66 ;
      RECT 6.24 203.46 8.21 204.26 ;
      RECT 6.24 200.06 8.21 200.86 ;
      RECT 6.24 196.66 8.21 197.46 ;
      RECT 6.24 193.26 8.21 194.06 ;
      RECT 6.24 189.86 8.21 190.66 ;
      RECT 6.24 186.46 8.21 187.26 ;
      RECT 6.24 183.06 8.21 183.86 ;
      RECT 6.24 179.66 8.21 180.46 ;
      RECT 6.24 176.26 8.21 177.06 ;
      RECT 6.24 172.86 8.21 173.66 ;
      RECT 6.24 169.46 8.21 170.26 ;
      RECT 6.24 166.06 8.21 166.86 ;
      RECT 6.24 162.66 8.21 163.46 ;
      RECT 6.24 159.26 8.21 160.06 ;
      RECT 6.24 155.86 8.21 156.66 ;
      RECT 6.24 152.46 8.21 153.26 ;
      RECT 6.24 149.06 8.21 149.86 ;
      RECT 6.24 145.66 8.21 146.46 ;
      RECT 6.24 142.26 8.21 143.06 ;
      RECT 6.24 138.86 8.21 139.66 ;
      RECT 6.24 135.46 8.21 136.26 ;
      RECT 6.24 132.06 8.21 132.86 ;
      RECT 6.24 128.66 8.21 129.46 ;
      RECT 6.24 125.26 8.21 126.06 ;
      RECT 6.24 121.86 8.21 122.66 ;
      RECT 6.24 118.46 8.21 119.26 ;
      RECT 6.24 115.06 8.21 115.86 ;
      RECT 6.24 111.66 8.21 112.46 ;
      RECT 6.24 108.26 8.21 109.06 ;
      RECT 6.24 104.86 8.21 105.66 ;
      RECT 6.24 101.46 8.21 102.26 ;
      RECT 6.24 98.06 8.21 98.86 ;
      RECT 6.24 94.66 8.21 95.46 ;
      RECT 6.24 91.26 8.21 92.06 ;
      RECT 6.24 87.86 8.21 88.66 ;
      RECT 6.24 84.46 8.21 85.26 ;
      RECT 6.24 81.06 8.21 81.86 ;
      RECT 6.24 77.66 8.21 78.46 ;
      RECT 6.24 74.26 8.21 75.06 ;
      RECT 6.24 70.86 8.21 71.66 ;
      RECT 7.41 3.12 9.41 67.05 ;
      RECT 6.24 54.22 9.41 55.22 ;
      RECT 6.24 41.29 9.41 42.29 ;
      RECT 6.24 39.44 9.41 40.44 ;
      RECT 6.24 32.98 9.41 33.98 ;
      RECT 6.24 31.13 9.41 32.13 ;
      RECT 6.24 21.41 9.41 22.21 ;
      RECT 6.24 12.64 9.41 13.74 ;
      RECT 6.24 505.6 6.84 506 ;
      RECT 6.44 504.36 6.84 506 ;
      RECT 6.24 504.36 6.84 505.16 ;
      RECT 238.6 0 240.6 517.18 ;
      RECT 235.48 3.12 237.48 514.06 ;
      RECT 233.76 7.94 234.36 9.14 ;
      RECT 233.76 17.26 234.36 18.46 ;
      RECT 233.76 25.81 234.36 27.81 ;
      RECT 233.76 35.91 234.36 36.91 ;
      RECT 233.76 50.24 234.36 51.24 ;
      RECT 233.76 57.02 234.36 58.02 ;
      RECT 233.76 60.6 234.36 61.6 ;
      RECT 233.76 62.45 234.36 63.45 ;
      RECT 233.76 69.16 234.36 69.96 ;
      RECT 233.76 72.56 234.36 73.36 ;
      RECT 233.76 75.96 234.36 76.76 ;
      RECT 233.76 79.36 234.36 80.16 ;
      RECT 233.76 82.76 234.36 83.56 ;
      RECT 233.76 86.16 234.36 86.96 ;
      RECT 233.76 89.56 234.36 90.36 ;
      RECT 233.76 92.96 234.36 93.76 ;
      RECT 233.76 96.36 234.36 97.16 ;
      RECT 233.76 99.76 234.36 100.56 ;
      RECT 233.76 103.16 234.36 103.96 ;
      RECT 233.76 106.56 234.36 107.36 ;
      RECT 233.76 109.96 234.36 110.76 ;
      RECT 233.76 113.36 234.36 114.16 ;
      RECT 233.76 116.76 234.36 117.56 ;
      RECT 233.76 120.16 234.36 120.96 ;
      RECT 233.76 123.56 234.36 124.36 ;
      RECT 233.76 126.96 234.36 127.76 ;
      RECT 233.76 130.36 234.36 131.16 ;
      RECT 233.76 133.76 234.36 134.56 ;
      RECT 233.76 137.16 234.36 137.96 ;
      RECT 233.76 140.56 234.36 141.36 ;
      RECT 233.76 143.96 234.36 144.76 ;
      RECT 233.76 147.36 234.36 148.16 ;
      RECT 233.76 150.76 234.36 151.56 ;
      RECT 233.76 154.16 234.36 154.96 ;
      RECT 233.76 157.56 234.36 158.36 ;
      RECT 233.76 160.96 234.36 161.76 ;
      RECT 233.76 164.36 234.36 165.16 ;
      RECT 233.76 167.76 234.36 168.56 ;
      RECT 233.76 171.16 234.36 171.96 ;
      RECT 233.76 174.56 234.36 175.36 ;
      RECT 233.76 177.96 234.36 178.76 ;
      RECT 233.76 181.36 234.36 182.16 ;
      RECT 233.76 184.76 234.36 185.56 ;
      RECT 233.76 188.16 234.36 188.96 ;
      RECT 233.76 191.56 234.36 192.36 ;
      RECT 233.76 194.96 234.36 195.76 ;
      RECT 233.76 198.36 234.36 199.16 ;
      RECT 233.76 201.76 234.36 202.56 ;
      RECT 233.76 205.16 234.36 205.96 ;
      RECT 233.76 208.56 234.36 209.36 ;
      RECT 233.76 211.96 234.36 212.76 ;
      RECT 233.76 215.36 234.36 216.16 ;
      RECT 233.76 218.76 234.36 219.56 ;
      RECT 233.76 222.16 234.36 222.96 ;
      RECT 233.76 225.56 234.36 226.36 ;
      RECT 233.76 228.96 234.36 229.76 ;
      RECT 233.76 232.36 234.36 233.16 ;
      RECT 233.76 235.76 234.36 236.56 ;
      RECT 233.76 239.16 234.36 239.96 ;
      RECT 233.76 242.56 234.36 243.36 ;
      RECT 233.76 245.96 234.36 246.76 ;
      RECT 233.76 249.36 234.36 250.16 ;
      RECT 233.76 252.76 234.36 253.56 ;
      RECT 233.76 256.16 234.36 256.96 ;
      RECT 233.76 259.56 234.36 260.36 ;
      RECT 233.76 262.96 234.36 263.76 ;
      RECT 233.76 266.36 234.36 267.16 ;
      RECT 233.76 269.76 234.36 270.56 ;
      RECT 233.76 273.16 234.36 273.96 ;
      RECT 233.76 276.56 234.36 277.36 ;
      RECT 233.76 279.96 234.36 280.76 ;
      RECT 233.76 283.36 234.36 284.16 ;
      RECT 233.76 286.76 234.36 287.56 ;
      RECT 233.76 290.16 234.36 290.96 ;
      RECT 233.76 293.56 234.36 294.36 ;
      RECT 233.76 296.96 234.36 297.76 ;
      RECT 233.76 300.36 234.36 301.16 ;
      RECT 233.76 303.76 234.36 304.56 ;
      RECT 233.76 307.16 234.36 307.96 ;
      RECT 233.76 310.56 234.36 311.36 ;
      RECT 233.76 313.96 234.36 314.76 ;
      RECT 233.76 317.36 234.36 318.16 ;
      RECT 233.76 320.76 234.36 321.56 ;
      RECT 233.76 324.16 234.36 324.96 ;
      RECT 233.76 327.56 234.36 328.36 ;
      RECT 233.76 330.96 234.36 331.76 ;
      RECT 233.76 334.36 234.36 335.16 ;
      RECT 233.76 337.76 234.36 338.56 ;
      RECT 233.76 341.16 234.36 341.96 ;
      RECT 233.76 344.56 234.36 345.36 ;
      RECT 233.76 347.96 234.36 348.76 ;
      RECT 233.76 351.36 234.36 352.16 ;
      RECT 233.76 354.76 234.36 355.56 ;
      RECT 233.76 358.16 234.36 358.96 ;
      RECT 233.76 361.56 234.36 362.36 ;
      RECT 233.76 364.96 234.36 365.76 ;
      RECT 233.76 368.36 234.36 369.16 ;
      RECT 233.76 371.76 234.36 372.56 ;
      RECT 233.76 375.16 234.36 375.96 ;
      RECT 233.76 378.56 234.36 379.36 ;
      RECT 233.76 381.96 234.36 382.76 ;
      RECT 233.76 385.36 234.36 386.16 ;
      RECT 233.76 388.76 234.36 389.56 ;
      RECT 233.76 392.16 234.36 392.96 ;
      RECT 233.76 395.56 234.36 396.36 ;
      RECT 233.76 398.96 234.36 399.76 ;
      RECT 233.76 402.36 234.36 403.16 ;
      RECT 233.76 405.76 234.36 406.56 ;
      RECT 233.76 409.16 234.36 409.96 ;
      RECT 233.76 412.56 234.36 413.36 ;
      RECT 233.76 415.96 234.36 416.76 ;
      RECT 233.76 419.36 234.36 420.16 ;
      RECT 233.76 422.76 234.36 423.56 ;
      RECT 233.76 426.16 234.36 426.96 ;
      RECT 233.76 429.56 234.36 430.36 ;
      RECT 233.76 432.96 234.36 433.76 ;
      RECT 233.76 436.36 234.36 437.16 ;
      RECT 233.76 439.76 234.36 440.56 ;
      RECT 233.76 443.16 234.36 443.96 ;
      RECT 233.76 446.56 234.36 447.36 ;
      RECT 233.76 449.96 234.36 450.76 ;
      RECT 233.76 453.36 234.36 454.16 ;
      RECT 233.76 456.76 234.36 457.56 ;
      RECT 233.76 460.16 234.36 460.96 ;
      RECT 233.76 463.56 234.36 464.36 ;
      RECT 233.76 466.96 234.36 467.76 ;
      RECT 233.76 470.36 234.36 471.16 ;
      RECT 233.76 473.76 234.36 474.56 ;
      RECT 233.76 477.16 234.36 477.96 ;
      RECT 233.76 480.56 234.36 481.36 ;
      RECT 233.76 483.96 234.36 484.76 ;
      RECT 233.76 487.36 234.36 488.16 ;
      RECT 233.76 490.76 234.36 491.56 ;
      RECT 233.76 494.16 234.36 494.96 ;
      RECT 233.76 497.56 234.36 498.36 ;
      RECT 233.76 500.96 234.36 501.76 ;
      RECT 233.76 509 234.36 509.8 ;
      RECT 152.89 7.14 153.49 7.59 ;
      RECT 151.99 8.19 152.79 517.18 ;
      RECT 151.29 6.24 151.89 7.59 ;
      RECT 149.27 7.14 149.87 7.59 ;
      RECT 146.09 3.12 147.41 514.06 ;
      RECT 144.01 7.14 144.61 7.59 ;
      RECT 141.62 6.24 142.22 7.59 ;
      RECT 137.81 7.14 138.41 7.59 ;
      RECT 134.41 7.14 135.01 7.59 ;
      RECT 131.01 7.14 131.61 7.59 ;
      RECT 127.61 7.14 128.21 7.59 ;
      RECT 120.81 7.14 121.41 7.59 ;
      RECT 117.41 7.14 118.01 7.59 ;
      RECT 114.01 7.14 114.61 7.59 ;
      RECT 107.21 7.14 107.81 7.59 ;
      RECT 106.11 66.63 107.21 514.06 ;
      RECT 103.81 7.14 104.41 7.59 ;
      RECT 100.41 7.14 101.01 7.59 ;
      RECT 99.31 66.63 100.41 514.06 ;
      RECT 93.61 7.14 94.21 7.59 ;
      RECT 92.51 66.63 93.61 514.06 ;
      RECT 90.21 7.14 90.81 7.59 ;
      RECT 18.81 6.24 19.41 7.04 ;
      RECT 6.24 7.94 6.84 9.14 ;
      RECT 6.24 17.26 6.84 18.46 ;
      RECT 6.24 25.81 6.84 27.81 ;
      RECT 6.24 35.91 6.84 36.91 ;
      RECT 6.24 50.24 6.84 51.24 ;
      RECT 6.24 57.02 6.84 58.02 ;
      RECT 6.24 60.6 6.84 61.6 ;
      RECT 6.24 62.45 6.84 63.45 ;
      RECT 6.24 69.16 6.84 69.96 ;
      RECT 6.24 72.56 6.84 73.36 ;
      RECT 6.24 75.96 6.84 76.76 ;
      RECT 6.24 79.36 6.84 80.16 ;
      RECT 6.24 82.76 6.84 83.56 ;
      RECT 6.24 86.16 6.84 86.96 ;
      RECT 6.24 89.56 6.84 90.36 ;
      RECT 6.24 92.96 6.84 93.76 ;
      RECT 6.24 96.36 6.84 97.16 ;
      RECT 6.24 99.76 6.84 100.56 ;
      RECT 6.24 103.16 6.84 103.96 ;
      RECT 6.24 106.56 6.84 107.36 ;
      RECT 6.24 109.96 6.84 110.76 ;
      RECT 6.24 113.36 6.84 114.16 ;
      RECT 6.24 116.76 6.84 117.56 ;
      RECT 6.24 120.16 6.84 120.96 ;
      RECT 6.24 123.56 6.84 124.36 ;
      RECT 6.24 126.96 6.84 127.76 ;
      RECT 6.24 130.36 6.84 131.16 ;
      RECT 6.24 133.76 6.84 134.56 ;
      RECT 6.24 137.16 6.84 137.96 ;
      RECT 6.24 140.56 6.84 141.36 ;
      RECT 6.24 143.96 6.84 144.76 ;
      RECT 6.24 147.36 6.84 148.16 ;
      RECT 6.24 150.76 6.84 151.56 ;
      RECT 6.24 154.16 6.84 154.96 ;
      RECT 6.24 157.56 6.84 158.36 ;
      RECT 6.24 160.96 6.84 161.76 ;
      RECT 6.24 164.36 6.84 165.16 ;
      RECT 6.24 167.76 6.84 168.56 ;
      RECT 6.24 171.16 6.84 171.96 ;
      RECT 6.24 174.56 6.84 175.36 ;
      RECT 6.24 177.96 6.84 178.76 ;
      RECT 6.24 181.36 6.84 182.16 ;
      RECT 6.24 184.76 6.84 185.56 ;
      RECT 6.24 188.16 6.84 188.96 ;
      RECT 6.24 191.56 6.84 192.36 ;
      RECT 6.24 194.96 6.84 195.76 ;
      RECT 6.24 198.36 6.84 199.16 ;
      RECT 6.24 201.76 6.84 202.56 ;
      RECT 6.24 205.16 6.84 205.96 ;
      RECT 6.24 208.56 6.84 209.36 ;
      RECT 6.24 211.96 6.84 212.76 ;
      RECT 6.24 215.36 6.84 216.16 ;
      RECT 6.24 218.76 6.84 219.56 ;
      RECT 6.24 222.16 6.84 222.96 ;
      RECT 6.24 225.56 6.84 226.36 ;
      RECT 6.24 228.96 6.84 229.76 ;
      RECT 6.24 232.36 6.84 233.16 ;
      RECT 6.24 235.76 6.84 236.56 ;
      RECT 6.24 239.16 6.84 239.96 ;
      RECT 6.24 242.56 6.84 243.36 ;
      RECT 6.24 245.96 6.84 246.76 ;
      RECT 6.24 249.36 6.84 250.16 ;
      RECT 6.24 252.76 6.84 253.56 ;
      RECT 6.24 256.16 6.84 256.96 ;
      RECT 6.24 259.56 6.84 260.36 ;
      RECT 6.24 262.96 6.84 263.76 ;
      RECT 6.24 266.36 6.84 267.16 ;
      RECT 6.24 269.76 6.84 270.56 ;
      RECT 6.24 273.16 6.84 273.96 ;
      RECT 6.24 276.56 6.84 277.36 ;
      RECT 6.24 279.96 6.84 280.76 ;
      RECT 6.24 283.36 6.84 284.16 ;
      RECT 6.24 286.76 6.84 287.56 ;
      RECT 6.24 290.16 6.84 290.96 ;
      RECT 6.24 293.56 6.84 294.36 ;
      RECT 6.24 296.96 6.84 297.76 ;
      RECT 6.24 300.36 6.84 301.16 ;
      RECT 6.24 303.76 6.84 304.56 ;
      RECT 6.24 307.16 6.84 307.96 ;
      RECT 6.24 310.56 6.84 311.36 ;
      RECT 6.24 313.96 6.84 314.76 ;
      RECT 6.24 317.36 6.84 318.16 ;
      RECT 6.24 320.76 6.84 321.56 ;
      RECT 6.24 324.16 6.84 324.96 ;
      RECT 6.24 327.56 6.84 328.36 ;
      RECT 6.24 330.96 6.84 331.76 ;
      RECT 6.24 334.36 6.84 335.16 ;
      RECT 6.24 337.76 6.84 338.56 ;
      RECT 6.24 341.16 6.84 341.96 ;
      RECT 6.24 344.56 6.84 345.36 ;
      RECT 6.24 347.96 6.84 348.76 ;
      RECT 6.24 351.36 6.84 352.16 ;
      RECT 6.24 354.76 6.84 355.56 ;
      RECT 6.24 358.16 6.84 358.96 ;
      RECT 6.24 361.56 6.84 362.36 ;
      RECT 6.24 364.96 6.84 365.76 ;
      RECT 6.24 368.36 6.84 369.16 ;
      RECT 6.24 371.76 6.84 372.56 ;
      RECT 6.24 375.16 6.84 375.96 ;
      RECT 6.24 378.56 6.84 379.36 ;
      RECT 6.24 381.96 6.84 382.76 ;
      RECT 6.24 385.36 6.84 386.16 ;
      RECT 6.24 388.76 6.84 389.56 ;
      RECT 6.24 392.16 6.84 392.96 ;
      RECT 6.24 395.56 6.84 396.36 ;
      RECT 6.24 398.96 6.84 399.76 ;
      RECT 6.24 402.36 6.84 403.16 ;
      RECT 6.24 405.76 6.84 406.56 ;
      RECT 6.24 409.16 6.84 409.96 ;
      RECT 6.24 412.56 6.84 413.36 ;
      RECT 6.24 415.96 6.84 416.76 ;
      RECT 6.24 419.36 6.84 420.16 ;
      RECT 6.24 422.76 6.84 423.56 ;
      RECT 6.24 426.16 6.84 426.96 ;
      RECT 6.24 429.56 6.84 430.36 ;
      RECT 6.24 432.96 6.84 433.76 ;
      RECT 6.24 436.36 6.84 437.16 ;
      RECT 6.24 439.76 6.84 440.56 ;
      RECT 6.24 443.16 6.84 443.96 ;
      RECT 6.24 446.56 6.84 447.36 ;
      RECT 6.24 449.96 6.84 450.76 ;
      RECT 6.24 453.36 6.84 454.16 ;
      RECT 6.24 456.76 6.84 457.56 ;
      RECT 6.24 460.16 6.84 460.96 ;
      RECT 6.24 463.56 6.84 464.36 ;
      RECT 6.24 466.96 6.84 467.76 ;
      RECT 6.24 470.36 6.84 471.16 ;
      RECT 6.24 473.76 6.84 474.56 ;
      RECT 6.24 477.16 6.84 477.96 ;
      RECT 6.24 480.56 6.84 481.36 ;
      RECT 6.24 483.96 6.84 484.76 ;
      RECT 6.24 487.36 6.84 488.16 ;
      RECT 6.24 490.76 6.84 491.56 ;
      RECT 6.24 494.16 6.84 494.96 ;
      RECT 6.24 497.56 6.84 498.36 ;
      RECT 6.24 500.96 6.84 501.76 ;
      RECT 6.24 509 6.84 509.8 ;
      RECT 3.12 3.12 5.12 514.06 ;
      RECT 0 0 2 517.18 ;
  END
END RA1SHD

END LIBRARY
